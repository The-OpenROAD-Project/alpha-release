VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x95
  FOREIGN fakeram45_256x95 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 57.452 BY 167.760 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 166.220 0.140 166.360 ;
      LAYER metal2 ;
      RECT 0.000 166.220 0.140 166.360 ;
      LAYER metal3 ;
      RECT 0.000 166.220 0.140 166.360 ;
      LAYER metal4 ;
      RECT 0.000 166.220 0.140 166.360 ;
      END
    END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 165.663 0.140 165.803 ;
      LAYER metal2 ;
      RECT 0.000 165.663 0.140 165.803 ;
      LAYER metal3 ;
      RECT 0.000 165.663 0.140 165.803 ;
      LAYER metal4 ;
      RECT 0.000 165.663 0.140 165.803 ;
      END
    END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 165.106 0.140 165.246 ;
      LAYER metal2 ;
      RECT 0.000 165.106 0.140 165.246 ;
      LAYER metal3 ;
      RECT 0.000 165.106 0.140 165.246 ;
      LAYER metal4 ;
      RECT 0.000 165.106 0.140 165.246 ;
      END
    END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 164.548 0.140 164.688 ;
      LAYER metal2 ;
      RECT 0.000 164.548 0.140 164.688 ;
      LAYER metal3 ;
      RECT 0.000 164.548 0.140 164.688 ;
      LAYER metal4 ;
      RECT 0.000 164.548 0.140 164.688 ;
      END
    END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 163.991 0.140 164.131 ;
      LAYER metal2 ;
      RECT 0.000 163.991 0.140 164.131 ;
      LAYER metal3 ;
      RECT 0.000 163.991 0.140 164.131 ;
      LAYER metal4 ;
      RECT 0.000 163.991 0.140 164.131 ;
      END
    END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 163.434 0.140 163.574 ;
      LAYER metal2 ;
      RECT 0.000 163.434 0.140 163.574 ;
      LAYER metal3 ;
      RECT 0.000 163.434 0.140 163.574 ;
      LAYER metal4 ;
      RECT 0.000 163.434 0.140 163.574 ;
      END
    END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 162.876 0.140 163.016 ;
      LAYER metal2 ;
      RECT 0.000 162.876 0.140 163.016 ;
      LAYER metal3 ;
      RECT 0.000 162.876 0.140 163.016 ;
      LAYER metal4 ;
      RECT 0.000 162.876 0.140 163.016 ;
      END
    END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 162.319 0.140 162.459 ;
      LAYER metal2 ;
      RECT 0.000 162.319 0.140 162.459 ;
      LAYER metal3 ;
      RECT 0.000 162.319 0.140 162.459 ;
      LAYER metal4 ;
      RECT 0.000 162.319 0.140 162.459 ;
      END
    END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 161.762 0.140 161.902 ;
      LAYER metal2 ;
      RECT 0.000 161.762 0.140 161.902 ;
      LAYER metal3 ;
      RECT 0.000 161.762 0.140 161.902 ;
      LAYER metal4 ;
      RECT 0.000 161.762 0.140 161.902 ;
      END
    END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 161.204 0.140 161.344 ;
      LAYER metal2 ;
      RECT 0.000 161.204 0.140 161.344 ;
      LAYER metal3 ;
      RECT 0.000 161.204 0.140 161.344 ;
      LAYER metal4 ;
      RECT 0.000 161.204 0.140 161.344 ;
      END
    END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 160.647 0.140 160.787 ;
      LAYER metal2 ;
      RECT 0.000 160.647 0.140 160.787 ;
      LAYER metal3 ;
      RECT 0.000 160.647 0.140 160.787 ;
      LAYER metal4 ;
      RECT 0.000 160.647 0.140 160.787 ;
      END
    END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 160.090 0.140 160.230 ;
      LAYER metal2 ;
      RECT 0.000 160.090 0.140 160.230 ;
      LAYER metal3 ;
      RECT 0.000 160.090 0.140 160.230 ;
      LAYER metal4 ;
      RECT 0.000 160.090 0.140 160.230 ;
      END
    END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 159.533 0.140 159.673 ;
      LAYER metal2 ;
      RECT 0.000 159.533 0.140 159.673 ;
      LAYER metal3 ;
      RECT 0.000 159.533 0.140 159.673 ;
      LAYER metal4 ;
      RECT 0.000 159.533 0.140 159.673 ;
      END
    END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 158.975 0.140 159.115 ;
      LAYER metal2 ;
      RECT 0.000 158.975 0.140 159.115 ;
      LAYER metal3 ;
      RECT 0.000 158.975 0.140 159.115 ;
      LAYER metal4 ;
      RECT 0.000 158.975 0.140 159.115 ;
      END
    END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 158.418 0.140 158.558 ;
      LAYER metal2 ;
      RECT 0.000 158.418 0.140 158.558 ;
      LAYER metal3 ;
      RECT 0.000 158.418 0.140 158.558 ;
      LAYER metal4 ;
      RECT 0.000 158.418 0.140 158.558 ;
      END
    END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 157.861 0.140 158.001 ;
      LAYER metal2 ;
      RECT 0.000 157.861 0.140 158.001 ;
      LAYER metal3 ;
      RECT 0.000 157.861 0.140 158.001 ;
      LAYER metal4 ;
      RECT 0.000 157.861 0.140 158.001 ;
      END
    END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 157.303 0.140 157.443 ;
      LAYER metal2 ;
      RECT 0.000 157.303 0.140 157.443 ;
      LAYER metal3 ;
      RECT 0.000 157.303 0.140 157.443 ;
      LAYER metal4 ;
      RECT 0.000 157.303 0.140 157.443 ;
      END
    END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 156.746 0.140 156.886 ;
      LAYER metal2 ;
      RECT 0.000 156.746 0.140 156.886 ;
      LAYER metal3 ;
      RECT 0.000 156.746 0.140 156.886 ;
      LAYER metal4 ;
      RECT 0.000 156.746 0.140 156.886 ;
      END
    END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 156.189 0.140 156.329 ;
      LAYER metal2 ;
      RECT 0.000 156.189 0.140 156.329 ;
      LAYER metal3 ;
      RECT 0.000 156.189 0.140 156.329 ;
      LAYER metal4 ;
      RECT 0.000 156.189 0.140 156.329 ;
      END
    END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 155.631 0.140 155.771 ;
      LAYER metal2 ;
      RECT 0.000 155.631 0.140 155.771 ;
      LAYER metal3 ;
      RECT 0.000 155.631 0.140 155.771 ;
      LAYER metal4 ;
      RECT 0.000 155.631 0.140 155.771 ;
      END
    END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 155.074 0.140 155.214 ;
      LAYER metal2 ;
      RECT 0.000 155.074 0.140 155.214 ;
      LAYER metal3 ;
      RECT 0.000 155.074 0.140 155.214 ;
      LAYER metal4 ;
      RECT 0.000 155.074 0.140 155.214 ;
      END
    END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 154.517 0.140 154.657 ;
      LAYER metal2 ;
      RECT 0.000 154.517 0.140 154.657 ;
      LAYER metal3 ;
      RECT 0.000 154.517 0.140 154.657 ;
      LAYER metal4 ;
      RECT 0.000 154.517 0.140 154.657 ;
      END
    END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 153.960 0.140 154.100 ;
      LAYER metal2 ;
      RECT 0.000 153.960 0.140 154.100 ;
      LAYER metal3 ;
      RECT 0.000 153.960 0.140 154.100 ;
      LAYER metal4 ;
      RECT 0.000 153.960 0.140 154.100 ;
      END
    END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 153.402 0.140 153.542 ;
      LAYER metal2 ;
      RECT 0.000 153.402 0.140 153.542 ;
      LAYER metal3 ;
      RECT 0.000 153.402 0.140 153.542 ;
      LAYER metal4 ;
      RECT 0.000 153.402 0.140 153.542 ;
      END
    END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 152.845 0.140 152.985 ;
      LAYER metal2 ;
      RECT 0.000 152.845 0.140 152.985 ;
      LAYER metal3 ;
      RECT 0.000 152.845 0.140 152.985 ;
      LAYER metal4 ;
      RECT 0.000 152.845 0.140 152.985 ;
      END
    END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 152.288 0.140 152.428 ;
      LAYER metal2 ;
      RECT 0.000 152.288 0.140 152.428 ;
      LAYER metal3 ;
      RECT 0.000 152.288 0.140 152.428 ;
      LAYER metal4 ;
      RECT 0.000 152.288 0.140 152.428 ;
      END
    END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 151.730 0.140 151.870 ;
      LAYER metal2 ;
      RECT 0.000 151.730 0.140 151.870 ;
      LAYER metal3 ;
      RECT 0.000 151.730 0.140 151.870 ;
      LAYER metal4 ;
      RECT 0.000 151.730 0.140 151.870 ;
      END
    END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 151.173 0.140 151.313 ;
      LAYER metal2 ;
      RECT 0.000 151.173 0.140 151.313 ;
      LAYER metal3 ;
      RECT 0.000 151.173 0.140 151.313 ;
      LAYER metal4 ;
      RECT 0.000 151.173 0.140 151.313 ;
      END
    END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 150.616 0.140 150.756 ;
      LAYER metal2 ;
      RECT 0.000 150.616 0.140 150.756 ;
      LAYER metal3 ;
      RECT 0.000 150.616 0.140 150.756 ;
      LAYER metal4 ;
      RECT 0.000 150.616 0.140 150.756 ;
      END
    END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 150.059 0.140 150.199 ;
      LAYER metal2 ;
      RECT 0.000 150.059 0.140 150.199 ;
      LAYER metal3 ;
      RECT 0.000 150.059 0.140 150.199 ;
      LAYER metal4 ;
      RECT 0.000 150.059 0.140 150.199 ;
      END
    END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 149.501 0.140 149.641 ;
      LAYER metal2 ;
      RECT 0.000 149.501 0.140 149.641 ;
      LAYER metal3 ;
      RECT 0.000 149.501 0.140 149.641 ;
      LAYER metal4 ;
      RECT 0.000 149.501 0.140 149.641 ;
      END
    END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 148.944 0.140 149.084 ;
      LAYER metal2 ;
      RECT 0.000 148.944 0.140 149.084 ;
      LAYER metal3 ;
      RECT 0.000 148.944 0.140 149.084 ;
      LAYER metal4 ;
      RECT 0.000 148.944 0.140 149.084 ;
      END
    END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 148.387 0.140 148.527 ;
      LAYER metal2 ;
      RECT 0.000 148.387 0.140 148.527 ;
      LAYER metal3 ;
      RECT 0.000 148.387 0.140 148.527 ;
      LAYER metal4 ;
      RECT 0.000 148.387 0.140 148.527 ;
      END
    END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 147.829 0.140 147.969 ;
      LAYER metal2 ;
      RECT 0.000 147.829 0.140 147.969 ;
      LAYER metal3 ;
      RECT 0.000 147.829 0.140 147.969 ;
      LAYER metal4 ;
      RECT 0.000 147.829 0.140 147.969 ;
      END
    END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 147.272 0.140 147.412 ;
      LAYER metal2 ;
      RECT 0.000 147.272 0.140 147.412 ;
      LAYER metal3 ;
      RECT 0.000 147.272 0.140 147.412 ;
      LAYER metal4 ;
      RECT 0.000 147.272 0.140 147.412 ;
      END
    END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 146.715 0.140 146.855 ;
      LAYER metal2 ;
      RECT 0.000 146.715 0.140 146.855 ;
      LAYER metal3 ;
      RECT 0.000 146.715 0.140 146.855 ;
      LAYER metal4 ;
      RECT 0.000 146.715 0.140 146.855 ;
      END
    END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 146.157 0.140 146.297 ;
      LAYER metal2 ;
      RECT 0.000 146.157 0.140 146.297 ;
      LAYER metal3 ;
      RECT 0.000 146.157 0.140 146.297 ;
      LAYER metal4 ;
      RECT 0.000 146.157 0.140 146.297 ;
      END
    END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 145.600 0.140 145.740 ;
      LAYER metal2 ;
      RECT 0.000 145.600 0.140 145.740 ;
      LAYER metal3 ;
      RECT 0.000 145.600 0.140 145.740 ;
      LAYER metal4 ;
      RECT 0.000 145.600 0.140 145.740 ;
      END
    END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 145.043 0.140 145.183 ;
      LAYER metal2 ;
      RECT 0.000 145.043 0.140 145.183 ;
      LAYER metal3 ;
      RECT 0.000 145.043 0.140 145.183 ;
      LAYER metal4 ;
      RECT 0.000 145.043 0.140 145.183 ;
      END
    END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 144.486 0.140 144.626 ;
      LAYER metal2 ;
      RECT 0.000 144.486 0.140 144.626 ;
      LAYER metal3 ;
      RECT 0.000 144.486 0.140 144.626 ;
      LAYER metal4 ;
      RECT 0.000 144.486 0.140 144.626 ;
      END
    END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 143.928 0.140 144.068 ;
      LAYER metal2 ;
      RECT 0.000 143.928 0.140 144.068 ;
      LAYER metal3 ;
      RECT 0.000 143.928 0.140 144.068 ;
      LAYER metal4 ;
      RECT 0.000 143.928 0.140 144.068 ;
      END
    END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 143.371 0.140 143.511 ;
      LAYER metal2 ;
      RECT 0.000 143.371 0.140 143.511 ;
      LAYER metal3 ;
      RECT 0.000 143.371 0.140 143.511 ;
      LAYER metal4 ;
      RECT 0.000 143.371 0.140 143.511 ;
      END
    END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 142.814 0.140 142.954 ;
      LAYER metal2 ;
      RECT 0.000 142.814 0.140 142.954 ;
      LAYER metal3 ;
      RECT 0.000 142.814 0.140 142.954 ;
      LAYER metal4 ;
      RECT 0.000 142.814 0.140 142.954 ;
      END
    END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 142.256 0.140 142.396 ;
      LAYER metal2 ;
      RECT 0.000 142.256 0.140 142.396 ;
      LAYER metal3 ;
      RECT 0.000 142.256 0.140 142.396 ;
      LAYER metal4 ;
      RECT 0.000 142.256 0.140 142.396 ;
      END
    END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 141.699 0.140 141.839 ;
      LAYER metal2 ;
      RECT 0.000 141.699 0.140 141.839 ;
      LAYER metal3 ;
      RECT 0.000 141.699 0.140 141.839 ;
      LAYER metal4 ;
      RECT 0.000 141.699 0.140 141.839 ;
      END
    END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 141.142 0.140 141.282 ;
      LAYER metal2 ;
      RECT 0.000 141.142 0.140 141.282 ;
      LAYER metal3 ;
      RECT 0.000 141.142 0.140 141.282 ;
      LAYER metal4 ;
      RECT 0.000 141.142 0.140 141.282 ;
      END
    END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 140.584 0.140 140.724 ;
      LAYER metal2 ;
      RECT 0.000 140.584 0.140 140.724 ;
      LAYER metal3 ;
      RECT 0.000 140.584 0.140 140.724 ;
      LAYER metal4 ;
      RECT 0.000 140.584 0.140 140.724 ;
      END
    END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 140.027 0.140 140.167 ;
      LAYER metal2 ;
      RECT 0.000 140.027 0.140 140.167 ;
      LAYER metal3 ;
      RECT 0.000 140.027 0.140 140.167 ;
      LAYER metal4 ;
      RECT 0.000 140.027 0.140 140.167 ;
      END
    END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 139.470 0.140 139.610 ;
      LAYER metal2 ;
      RECT 0.000 139.470 0.140 139.610 ;
      LAYER metal3 ;
      RECT 0.000 139.470 0.140 139.610 ;
      LAYER metal4 ;
      RECT 0.000 139.470 0.140 139.610 ;
      END
    END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 138.913 0.140 139.053 ;
      LAYER metal2 ;
      RECT 0.000 138.913 0.140 139.053 ;
      LAYER metal3 ;
      RECT 0.000 138.913 0.140 139.053 ;
      LAYER metal4 ;
      RECT 0.000 138.913 0.140 139.053 ;
      END
    END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 138.355 0.140 138.495 ;
      LAYER metal2 ;
      RECT 0.000 138.355 0.140 138.495 ;
      LAYER metal3 ;
      RECT 0.000 138.355 0.140 138.495 ;
      LAYER metal4 ;
      RECT 0.000 138.355 0.140 138.495 ;
      END
    END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 137.798 0.140 137.938 ;
      LAYER metal2 ;
      RECT 0.000 137.798 0.140 137.938 ;
      LAYER metal3 ;
      RECT 0.000 137.798 0.140 137.938 ;
      LAYER metal4 ;
      RECT 0.000 137.798 0.140 137.938 ;
      END
    END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 137.241 0.140 137.381 ;
      LAYER metal2 ;
      RECT 0.000 137.241 0.140 137.381 ;
      LAYER metal3 ;
      RECT 0.000 137.241 0.140 137.381 ;
      LAYER metal4 ;
      RECT 0.000 137.241 0.140 137.381 ;
      END
    END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 136.683 0.140 136.823 ;
      LAYER metal2 ;
      RECT 0.000 136.683 0.140 136.823 ;
      LAYER metal3 ;
      RECT 0.000 136.683 0.140 136.823 ;
      LAYER metal4 ;
      RECT 0.000 136.683 0.140 136.823 ;
      END
    END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 136.126 0.140 136.266 ;
      LAYER metal2 ;
      RECT 0.000 136.126 0.140 136.266 ;
      LAYER metal3 ;
      RECT 0.000 136.126 0.140 136.266 ;
      LAYER metal4 ;
      RECT 0.000 136.126 0.140 136.266 ;
      END
    END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 135.569 0.140 135.709 ;
      LAYER metal2 ;
      RECT 0.000 135.569 0.140 135.709 ;
      LAYER metal3 ;
      RECT 0.000 135.569 0.140 135.709 ;
      LAYER metal4 ;
      RECT 0.000 135.569 0.140 135.709 ;
      END
    END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 135.011 0.140 135.151 ;
      LAYER metal2 ;
      RECT 0.000 135.011 0.140 135.151 ;
      LAYER metal3 ;
      RECT 0.000 135.011 0.140 135.151 ;
      LAYER metal4 ;
      RECT 0.000 135.011 0.140 135.151 ;
      END
    END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 134.454 0.140 134.594 ;
      LAYER metal2 ;
      RECT 0.000 134.454 0.140 134.594 ;
      LAYER metal3 ;
      RECT 0.000 134.454 0.140 134.594 ;
      LAYER metal4 ;
      RECT 0.000 134.454 0.140 134.594 ;
      END
    END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 133.897 0.140 134.037 ;
      LAYER metal2 ;
      RECT 0.000 133.897 0.140 134.037 ;
      LAYER metal3 ;
      RECT 0.000 133.897 0.140 134.037 ;
      LAYER metal4 ;
      RECT 0.000 133.897 0.140 134.037 ;
      END
    END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 133.340 0.140 133.480 ;
      LAYER metal2 ;
      RECT 0.000 133.340 0.140 133.480 ;
      LAYER metal3 ;
      RECT 0.000 133.340 0.140 133.480 ;
      LAYER metal4 ;
      RECT 0.000 133.340 0.140 133.480 ;
      END
    END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 132.782 0.140 132.922 ;
      LAYER metal2 ;
      RECT 0.000 132.782 0.140 132.922 ;
      LAYER metal3 ;
      RECT 0.000 132.782 0.140 132.922 ;
      LAYER metal4 ;
      RECT 0.000 132.782 0.140 132.922 ;
      END
    END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 132.225 0.140 132.365 ;
      LAYER metal2 ;
      RECT 0.000 132.225 0.140 132.365 ;
      LAYER metal3 ;
      RECT 0.000 132.225 0.140 132.365 ;
      LAYER metal4 ;
      RECT 0.000 132.225 0.140 132.365 ;
      END
    END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 131.668 0.140 131.808 ;
      LAYER metal2 ;
      RECT 0.000 131.668 0.140 131.808 ;
      LAYER metal3 ;
      RECT 0.000 131.668 0.140 131.808 ;
      LAYER metal4 ;
      RECT 0.000 131.668 0.140 131.808 ;
      END
    END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 131.110 0.140 131.250 ;
      LAYER metal2 ;
      RECT 0.000 131.110 0.140 131.250 ;
      LAYER metal3 ;
      RECT 0.000 131.110 0.140 131.250 ;
      LAYER metal4 ;
      RECT 0.000 131.110 0.140 131.250 ;
      END
    END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 130.553 0.140 130.693 ;
      LAYER metal2 ;
      RECT 0.000 130.553 0.140 130.693 ;
      LAYER metal3 ;
      RECT 0.000 130.553 0.140 130.693 ;
      LAYER metal4 ;
      RECT 0.000 130.553 0.140 130.693 ;
      END
    END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 129.996 0.140 130.136 ;
      LAYER metal2 ;
      RECT 0.000 129.996 0.140 130.136 ;
      LAYER metal3 ;
      RECT 0.000 129.996 0.140 130.136 ;
      LAYER metal4 ;
      RECT 0.000 129.996 0.140 130.136 ;
      END
    END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 129.438 0.140 129.578 ;
      LAYER metal2 ;
      RECT 0.000 129.438 0.140 129.578 ;
      LAYER metal3 ;
      RECT 0.000 129.438 0.140 129.578 ;
      LAYER metal4 ;
      RECT 0.000 129.438 0.140 129.578 ;
      END
    END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 128.881 0.140 129.021 ;
      LAYER metal2 ;
      RECT 0.000 128.881 0.140 129.021 ;
      LAYER metal3 ;
      RECT 0.000 128.881 0.140 129.021 ;
      LAYER metal4 ;
      RECT 0.000 128.881 0.140 129.021 ;
      END
    END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 128.324 0.140 128.464 ;
      LAYER metal2 ;
      RECT 0.000 128.324 0.140 128.464 ;
      LAYER metal3 ;
      RECT 0.000 128.324 0.140 128.464 ;
      LAYER metal4 ;
      RECT 0.000 128.324 0.140 128.464 ;
      END
    END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 127.767 0.140 127.907 ;
      LAYER metal2 ;
      RECT 0.000 127.767 0.140 127.907 ;
      LAYER metal3 ;
      RECT 0.000 127.767 0.140 127.907 ;
      LAYER metal4 ;
      RECT 0.000 127.767 0.140 127.907 ;
      END
    END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 127.209 0.140 127.349 ;
      LAYER metal2 ;
      RECT 0.000 127.209 0.140 127.349 ;
      LAYER metal3 ;
      RECT 0.000 127.209 0.140 127.349 ;
      LAYER metal4 ;
      RECT 0.000 127.209 0.140 127.349 ;
      END
    END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 126.652 0.140 126.792 ;
      LAYER metal2 ;
      RECT 0.000 126.652 0.140 126.792 ;
      LAYER metal3 ;
      RECT 0.000 126.652 0.140 126.792 ;
      LAYER metal4 ;
      RECT 0.000 126.652 0.140 126.792 ;
      END
    END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 126.095 0.140 126.235 ;
      LAYER metal2 ;
      RECT 0.000 126.095 0.140 126.235 ;
      LAYER metal3 ;
      RECT 0.000 126.095 0.140 126.235 ;
      LAYER metal4 ;
      RECT 0.000 126.095 0.140 126.235 ;
      END
    END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 125.537 0.140 125.677 ;
      LAYER metal2 ;
      RECT 0.000 125.537 0.140 125.677 ;
      LAYER metal3 ;
      RECT 0.000 125.537 0.140 125.677 ;
      LAYER metal4 ;
      RECT 0.000 125.537 0.140 125.677 ;
      END
    END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 124.980 0.140 125.120 ;
      LAYER metal2 ;
      RECT 0.000 124.980 0.140 125.120 ;
      LAYER metal3 ;
      RECT 0.000 124.980 0.140 125.120 ;
      LAYER metal4 ;
      RECT 0.000 124.980 0.140 125.120 ;
      END
    END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 124.423 0.140 124.563 ;
      LAYER metal2 ;
      RECT 0.000 124.423 0.140 124.563 ;
      LAYER metal3 ;
      RECT 0.000 124.423 0.140 124.563 ;
      LAYER metal4 ;
      RECT 0.000 124.423 0.140 124.563 ;
      END
    END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 123.866 0.140 124.006 ;
      LAYER metal2 ;
      RECT 0.000 123.866 0.140 124.006 ;
      LAYER metal3 ;
      RECT 0.000 123.866 0.140 124.006 ;
      LAYER metal4 ;
      RECT 0.000 123.866 0.140 124.006 ;
      END
    END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 123.308 0.140 123.448 ;
      LAYER metal2 ;
      RECT 0.000 123.308 0.140 123.448 ;
      LAYER metal3 ;
      RECT 0.000 123.308 0.140 123.448 ;
      LAYER metal4 ;
      RECT 0.000 123.308 0.140 123.448 ;
      END
    END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 122.751 0.140 122.891 ;
      LAYER metal2 ;
      RECT 0.000 122.751 0.140 122.891 ;
      LAYER metal3 ;
      RECT 0.000 122.751 0.140 122.891 ;
      LAYER metal4 ;
      RECT 0.000 122.751 0.140 122.891 ;
      END
    END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 122.194 0.140 122.334 ;
      LAYER metal2 ;
      RECT 0.000 122.194 0.140 122.334 ;
      LAYER metal3 ;
      RECT 0.000 122.194 0.140 122.334 ;
      LAYER metal4 ;
      RECT 0.000 122.194 0.140 122.334 ;
      END
    END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 121.636 0.140 121.776 ;
      LAYER metal2 ;
      RECT 0.000 121.636 0.140 121.776 ;
      LAYER metal3 ;
      RECT 0.000 121.636 0.140 121.776 ;
      LAYER metal4 ;
      RECT 0.000 121.636 0.140 121.776 ;
      END
    END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 121.079 0.140 121.219 ;
      LAYER metal2 ;
      RECT 0.000 121.079 0.140 121.219 ;
      LAYER metal3 ;
      RECT 0.000 121.079 0.140 121.219 ;
      LAYER metal4 ;
      RECT 0.000 121.079 0.140 121.219 ;
      END
    END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 120.522 0.140 120.662 ;
      LAYER metal2 ;
      RECT 0.000 120.522 0.140 120.662 ;
      LAYER metal3 ;
      RECT 0.000 120.522 0.140 120.662 ;
      LAYER metal4 ;
      RECT 0.000 120.522 0.140 120.662 ;
      END
    END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 119.964 0.140 120.104 ;
      LAYER metal2 ;
      RECT 0.000 119.964 0.140 120.104 ;
      LAYER metal3 ;
      RECT 0.000 119.964 0.140 120.104 ;
      LAYER metal4 ;
      RECT 0.000 119.964 0.140 120.104 ;
      END
    END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 119.407 0.140 119.547 ;
      LAYER metal2 ;
      RECT 0.000 119.407 0.140 119.547 ;
      LAYER metal3 ;
      RECT 0.000 119.407 0.140 119.547 ;
      LAYER metal4 ;
      RECT 0.000 119.407 0.140 119.547 ;
      END
    END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 118.850 0.140 118.990 ;
      LAYER metal2 ;
      RECT 0.000 118.850 0.140 118.990 ;
      LAYER metal3 ;
      RECT 0.000 118.850 0.140 118.990 ;
      LAYER metal4 ;
      RECT 0.000 118.850 0.140 118.990 ;
      END
    END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 118.293 0.140 118.433 ;
      LAYER metal2 ;
      RECT 0.000 118.293 0.140 118.433 ;
      LAYER metal3 ;
      RECT 0.000 118.293 0.140 118.433 ;
      LAYER metal4 ;
      RECT 0.000 118.293 0.140 118.433 ;
      END
    END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 117.735 0.140 117.875 ;
      LAYER metal2 ;
      RECT 0.000 117.735 0.140 117.875 ;
      LAYER metal3 ;
      RECT 0.000 117.735 0.140 117.875 ;
      LAYER metal4 ;
      RECT 0.000 117.735 0.140 117.875 ;
      END
    END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 117.178 0.140 117.318 ;
      LAYER metal2 ;
      RECT 0.000 117.178 0.140 117.318 ;
      LAYER metal3 ;
      RECT 0.000 117.178 0.140 117.318 ;
      LAYER metal4 ;
      RECT 0.000 117.178 0.140 117.318 ;
      END
    END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 116.621 0.140 116.761 ;
      LAYER metal2 ;
      RECT 0.000 116.621 0.140 116.761 ;
      LAYER metal3 ;
      RECT 0.000 116.621 0.140 116.761 ;
      LAYER metal4 ;
      RECT 0.000 116.621 0.140 116.761 ;
      END
    END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 116.063 0.140 116.203 ;
      LAYER metal2 ;
      RECT 0.000 116.063 0.140 116.203 ;
      LAYER metal3 ;
      RECT 0.000 116.063 0.140 116.203 ;
      LAYER metal4 ;
      RECT 0.000 116.063 0.140 116.203 ;
      END
    END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 115.506 0.140 115.646 ;
      LAYER metal2 ;
      RECT 0.000 115.506 0.140 115.646 ;
      LAYER metal3 ;
      RECT 0.000 115.506 0.140 115.646 ;
      LAYER metal4 ;
      RECT 0.000 115.506 0.140 115.646 ;
      END
    END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 114.949 0.140 115.089 ;
      LAYER metal2 ;
      RECT 0.000 114.949 0.140 115.089 ;
      LAYER metal3 ;
      RECT 0.000 114.949 0.140 115.089 ;
      LAYER metal4 ;
      RECT 0.000 114.949 0.140 115.089 ;
      END
    END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 114.391 0.140 114.531 ;
      LAYER metal2 ;
      RECT 0.000 114.391 0.140 114.531 ;
      LAYER metal3 ;
      RECT 0.000 114.391 0.140 114.531 ;
      LAYER metal4 ;
      RECT 0.000 114.391 0.140 114.531 ;
      END
    END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 113.834 0.140 113.974 ;
      LAYER metal2 ;
      RECT 0.000 113.834 0.140 113.974 ;
      LAYER metal3 ;
      RECT 0.000 113.834 0.140 113.974 ;
      LAYER metal4 ;
      RECT 0.000 113.834 0.140 113.974 ;
      END
    END w_mask_in[94]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 113.277 0.140 113.417 ;
      LAYER metal2 ;
      RECT 0.000 113.277 0.140 113.417 ;
      LAYER metal3 ;
      RECT 0.000 113.277 0.140 113.417 ;
      LAYER metal4 ;
      RECT 0.000 113.277 0.140 113.417 ;
      END
    END we_in
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 112.720 0.140 112.860 ;
      LAYER metal2 ;
      RECT 0.000 112.720 0.140 112.860 ;
      LAYER metal3 ;
      RECT 0.000 112.720 0.140 112.860 ;
      LAYER metal4 ;
      RECT 0.000 112.720 0.140 112.860 ;
      END
    END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 112.162 0.140 112.302 ;
      LAYER metal2 ;
      RECT 0.000 112.162 0.140 112.302 ;
      LAYER metal3 ;
      RECT 0.000 112.162 0.140 112.302 ;
      LAYER metal4 ;
      RECT 0.000 112.162 0.140 112.302 ;
      END
    END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 111.605 0.140 111.745 ;
      LAYER metal2 ;
      RECT 0.000 111.605 0.140 111.745 ;
      LAYER metal3 ;
      RECT 0.000 111.605 0.140 111.745 ;
      LAYER metal4 ;
      RECT 0.000 111.605 0.140 111.745 ;
      END
    END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 111.048 0.140 111.188 ;
      LAYER metal2 ;
      RECT 0.000 111.048 0.140 111.188 ;
      LAYER metal3 ;
      RECT 0.000 111.048 0.140 111.188 ;
      LAYER metal4 ;
      RECT 0.000 111.048 0.140 111.188 ;
      END
    END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 110.490 0.140 110.630 ;
      LAYER metal2 ;
      RECT 0.000 110.490 0.140 110.630 ;
      LAYER metal3 ;
      RECT 0.000 110.490 0.140 110.630 ;
      LAYER metal4 ;
      RECT 0.000 110.490 0.140 110.630 ;
      END
    END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 109.933 0.140 110.073 ;
      LAYER metal2 ;
      RECT 0.000 109.933 0.140 110.073 ;
      LAYER metal3 ;
      RECT 0.000 109.933 0.140 110.073 ;
      LAYER metal4 ;
      RECT 0.000 109.933 0.140 110.073 ;
      END
    END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 109.376 0.140 109.516 ;
      LAYER metal2 ;
      RECT 0.000 109.376 0.140 109.516 ;
      LAYER metal3 ;
      RECT 0.000 109.376 0.140 109.516 ;
      LAYER metal4 ;
      RECT 0.000 109.376 0.140 109.516 ;
      END
    END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 108.818 0.140 108.958 ;
      LAYER metal2 ;
      RECT 0.000 108.818 0.140 108.958 ;
      LAYER metal3 ;
      RECT 0.000 108.818 0.140 108.958 ;
      LAYER metal4 ;
      RECT 0.000 108.818 0.140 108.958 ;
      END
    END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 108.261 0.140 108.401 ;
      LAYER metal2 ;
      RECT 0.000 108.261 0.140 108.401 ;
      LAYER metal3 ;
      RECT 0.000 108.261 0.140 108.401 ;
      LAYER metal4 ;
      RECT 0.000 108.261 0.140 108.401 ;
      END
    END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 107.704 0.140 107.844 ;
      LAYER metal2 ;
      RECT 0.000 107.704 0.140 107.844 ;
      LAYER metal3 ;
      RECT 0.000 107.704 0.140 107.844 ;
      LAYER metal4 ;
      RECT 0.000 107.704 0.140 107.844 ;
      END
    END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 107.147 0.140 107.287 ;
      LAYER metal2 ;
      RECT 0.000 107.147 0.140 107.287 ;
      LAYER metal3 ;
      RECT 0.000 107.147 0.140 107.287 ;
      LAYER metal4 ;
      RECT 0.000 107.147 0.140 107.287 ;
      END
    END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 106.589 0.140 106.729 ;
      LAYER metal2 ;
      RECT 0.000 106.589 0.140 106.729 ;
      LAYER metal3 ;
      RECT 0.000 106.589 0.140 106.729 ;
      LAYER metal4 ;
      RECT 0.000 106.589 0.140 106.729 ;
      END
    END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 106.032 0.140 106.172 ;
      LAYER metal2 ;
      RECT 0.000 106.032 0.140 106.172 ;
      LAYER metal3 ;
      RECT 0.000 106.032 0.140 106.172 ;
      LAYER metal4 ;
      RECT 0.000 106.032 0.140 106.172 ;
      END
    END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 105.475 0.140 105.615 ;
      LAYER metal2 ;
      RECT 0.000 105.475 0.140 105.615 ;
      LAYER metal3 ;
      RECT 0.000 105.475 0.140 105.615 ;
      LAYER metal4 ;
      RECT 0.000 105.475 0.140 105.615 ;
      END
    END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 104.917 0.140 105.057 ;
      LAYER metal2 ;
      RECT 0.000 104.917 0.140 105.057 ;
      LAYER metal3 ;
      RECT 0.000 104.917 0.140 105.057 ;
      LAYER metal4 ;
      RECT 0.000 104.917 0.140 105.057 ;
      END
    END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 104.360 0.140 104.500 ;
      LAYER metal2 ;
      RECT 0.000 104.360 0.140 104.500 ;
      LAYER metal3 ;
      RECT 0.000 104.360 0.140 104.500 ;
      LAYER metal4 ;
      RECT 0.000 104.360 0.140 104.500 ;
      END
    END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 103.803 0.140 103.943 ;
      LAYER metal2 ;
      RECT 0.000 103.803 0.140 103.943 ;
      LAYER metal3 ;
      RECT 0.000 103.803 0.140 103.943 ;
      LAYER metal4 ;
      RECT 0.000 103.803 0.140 103.943 ;
      END
    END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 103.245 0.140 103.385 ;
      LAYER metal2 ;
      RECT 0.000 103.245 0.140 103.385 ;
      LAYER metal3 ;
      RECT 0.000 103.245 0.140 103.385 ;
      LAYER metal4 ;
      RECT 0.000 103.245 0.140 103.385 ;
      END
    END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 102.688 0.140 102.828 ;
      LAYER metal2 ;
      RECT 0.000 102.688 0.140 102.828 ;
      LAYER metal3 ;
      RECT 0.000 102.688 0.140 102.828 ;
      LAYER metal4 ;
      RECT 0.000 102.688 0.140 102.828 ;
      END
    END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 102.131 0.140 102.271 ;
      LAYER metal2 ;
      RECT 0.000 102.131 0.140 102.271 ;
      LAYER metal3 ;
      RECT 0.000 102.131 0.140 102.271 ;
      LAYER metal4 ;
      RECT 0.000 102.131 0.140 102.271 ;
      END
    END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 101.574 0.140 101.714 ;
      LAYER metal2 ;
      RECT 0.000 101.574 0.140 101.714 ;
      LAYER metal3 ;
      RECT 0.000 101.574 0.140 101.714 ;
      LAYER metal4 ;
      RECT 0.000 101.574 0.140 101.714 ;
      END
    END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 101.016 0.140 101.156 ;
      LAYER metal2 ;
      RECT 0.000 101.016 0.140 101.156 ;
      LAYER metal3 ;
      RECT 0.000 101.016 0.140 101.156 ;
      LAYER metal4 ;
      RECT 0.000 101.016 0.140 101.156 ;
      END
    END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 100.459 0.140 100.599 ;
      LAYER metal2 ;
      RECT 0.000 100.459 0.140 100.599 ;
      LAYER metal3 ;
      RECT 0.000 100.459 0.140 100.599 ;
      LAYER metal4 ;
      RECT 0.000 100.459 0.140 100.599 ;
      END
    END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 99.902 0.140 100.042 ;
      LAYER metal2 ;
      RECT 0.000 99.902 0.140 100.042 ;
      LAYER metal3 ;
      RECT 0.000 99.902 0.140 100.042 ;
      LAYER metal4 ;
      RECT 0.000 99.902 0.140 100.042 ;
      END
    END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 99.344 0.140 99.484 ;
      LAYER metal2 ;
      RECT 0.000 99.344 0.140 99.484 ;
      LAYER metal3 ;
      RECT 0.000 99.344 0.140 99.484 ;
      LAYER metal4 ;
      RECT 0.000 99.344 0.140 99.484 ;
      END
    END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 98.787 0.140 98.927 ;
      LAYER metal2 ;
      RECT 0.000 98.787 0.140 98.927 ;
      LAYER metal3 ;
      RECT 0.000 98.787 0.140 98.927 ;
      LAYER metal4 ;
      RECT 0.000 98.787 0.140 98.927 ;
      END
    END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 98.230 0.140 98.370 ;
      LAYER metal2 ;
      RECT 0.000 98.230 0.140 98.370 ;
      LAYER metal3 ;
      RECT 0.000 98.230 0.140 98.370 ;
      LAYER metal4 ;
      RECT 0.000 98.230 0.140 98.370 ;
      END
    END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 97.673 0.140 97.813 ;
      LAYER metal2 ;
      RECT 0.000 97.673 0.140 97.813 ;
      LAYER metal3 ;
      RECT 0.000 97.673 0.140 97.813 ;
      LAYER metal4 ;
      RECT 0.000 97.673 0.140 97.813 ;
      END
    END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 97.115 0.140 97.255 ;
      LAYER metal2 ;
      RECT 0.000 97.115 0.140 97.255 ;
      LAYER metal3 ;
      RECT 0.000 97.115 0.140 97.255 ;
      LAYER metal4 ;
      RECT 0.000 97.115 0.140 97.255 ;
      END
    END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 96.558 0.140 96.698 ;
      LAYER metal2 ;
      RECT 0.000 96.558 0.140 96.698 ;
      LAYER metal3 ;
      RECT 0.000 96.558 0.140 96.698 ;
      LAYER metal4 ;
      RECT 0.000 96.558 0.140 96.698 ;
      END
    END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 96.001 0.140 96.141 ;
      LAYER metal2 ;
      RECT 0.000 96.001 0.140 96.141 ;
      LAYER metal3 ;
      RECT 0.000 96.001 0.140 96.141 ;
      LAYER metal4 ;
      RECT 0.000 96.001 0.140 96.141 ;
      END
    END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 95.443 0.140 95.583 ;
      LAYER metal2 ;
      RECT 0.000 95.443 0.140 95.583 ;
      LAYER metal3 ;
      RECT 0.000 95.443 0.140 95.583 ;
      LAYER metal4 ;
      RECT 0.000 95.443 0.140 95.583 ;
      END
    END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 94.886 0.140 95.026 ;
      LAYER metal2 ;
      RECT 0.000 94.886 0.140 95.026 ;
      LAYER metal3 ;
      RECT 0.000 94.886 0.140 95.026 ;
      LAYER metal4 ;
      RECT 0.000 94.886 0.140 95.026 ;
      END
    END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 94.329 0.140 94.469 ;
      LAYER metal2 ;
      RECT 0.000 94.329 0.140 94.469 ;
      LAYER metal3 ;
      RECT 0.000 94.329 0.140 94.469 ;
      LAYER metal4 ;
      RECT 0.000 94.329 0.140 94.469 ;
      END
    END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 93.771 0.140 93.911 ;
      LAYER metal2 ;
      RECT 0.000 93.771 0.140 93.911 ;
      LAYER metal3 ;
      RECT 0.000 93.771 0.140 93.911 ;
      LAYER metal4 ;
      RECT 0.000 93.771 0.140 93.911 ;
      END
    END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 93.214 0.140 93.354 ;
      LAYER metal2 ;
      RECT 0.000 93.214 0.140 93.354 ;
      LAYER metal3 ;
      RECT 0.000 93.214 0.140 93.354 ;
      LAYER metal4 ;
      RECT 0.000 93.214 0.140 93.354 ;
      END
    END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 92.657 0.140 92.797 ;
      LAYER metal2 ;
      RECT 0.000 92.657 0.140 92.797 ;
      LAYER metal3 ;
      RECT 0.000 92.657 0.140 92.797 ;
      LAYER metal4 ;
      RECT 0.000 92.657 0.140 92.797 ;
      END
    END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 92.100 0.140 92.240 ;
      LAYER metal2 ;
      RECT 0.000 92.100 0.140 92.240 ;
      LAYER metal3 ;
      RECT 0.000 92.100 0.140 92.240 ;
      LAYER metal4 ;
      RECT 0.000 92.100 0.140 92.240 ;
      END
    END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 91.542 0.140 91.682 ;
      LAYER metal2 ;
      RECT 0.000 91.542 0.140 91.682 ;
      LAYER metal3 ;
      RECT 0.000 91.542 0.140 91.682 ;
      LAYER metal4 ;
      RECT 0.000 91.542 0.140 91.682 ;
      END
    END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 90.985 0.140 91.125 ;
      LAYER metal2 ;
      RECT 0.000 90.985 0.140 91.125 ;
      LAYER metal3 ;
      RECT 0.000 90.985 0.140 91.125 ;
      LAYER metal4 ;
      RECT 0.000 90.985 0.140 91.125 ;
      END
    END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 90.428 0.140 90.568 ;
      LAYER metal2 ;
      RECT 0.000 90.428 0.140 90.568 ;
      LAYER metal3 ;
      RECT 0.000 90.428 0.140 90.568 ;
      LAYER metal4 ;
      RECT 0.000 90.428 0.140 90.568 ;
      END
    END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 89.870 0.140 90.010 ;
      LAYER metal2 ;
      RECT 0.000 89.870 0.140 90.010 ;
      LAYER metal3 ;
      RECT 0.000 89.870 0.140 90.010 ;
      LAYER metal4 ;
      RECT 0.000 89.870 0.140 90.010 ;
      END
    END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 89.313 0.140 89.453 ;
      LAYER metal2 ;
      RECT 0.000 89.313 0.140 89.453 ;
      LAYER metal3 ;
      RECT 0.000 89.313 0.140 89.453 ;
      LAYER metal4 ;
      RECT 0.000 89.313 0.140 89.453 ;
      END
    END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 88.756 0.140 88.896 ;
      LAYER metal2 ;
      RECT 0.000 88.756 0.140 88.896 ;
      LAYER metal3 ;
      RECT 0.000 88.756 0.140 88.896 ;
      LAYER metal4 ;
      RECT 0.000 88.756 0.140 88.896 ;
      END
    END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 88.198 0.140 88.338 ;
      LAYER metal2 ;
      RECT 0.000 88.198 0.140 88.338 ;
      LAYER metal3 ;
      RECT 0.000 88.198 0.140 88.338 ;
      LAYER metal4 ;
      RECT 0.000 88.198 0.140 88.338 ;
      END
    END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 87.641 0.140 87.781 ;
      LAYER metal2 ;
      RECT 0.000 87.641 0.140 87.781 ;
      LAYER metal3 ;
      RECT 0.000 87.641 0.140 87.781 ;
      LAYER metal4 ;
      RECT 0.000 87.641 0.140 87.781 ;
      END
    END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 87.084 0.140 87.224 ;
      LAYER metal2 ;
      RECT 0.000 87.084 0.140 87.224 ;
      LAYER metal3 ;
      RECT 0.000 87.084 0.140 87.224 ;
      LAYER metal4 ;
      RECT 0.000 87.084 0.140 87.224 ;
      END
    END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 86.527 0.140 86.667 ;
      LAYER metal2 ;
      RECT 0.000 86.527 0.140 86.667 ;
      LAYER metal3 ;
      RECT 0.000 86.527 0.140 86.667 ;
      LAYER metal4 ;
      RECT 0.000 86.527 0.140 86.667 ;
      END
    END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 85.969 0.140 86.109 ;
      LAYER metal2 ;
      RECT 0.000 85.969 0.140 86.109 ;
      LAYER metal3 ;
      RECT 0.000 85.969 0.140 86.109 ;
      LAYER metal4 ;
      RECT 0.000 85.969 0.140 86.109 ;
      END
    END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 85.412 0.140 85.552 ;
      LAYER metal2 ;
      RECT 0.000 85.412 0.140 85.552 ;
      LAYER metal3 ;
      RECT 0.000 85.412 0.140 85.552 ;
      LAYER metal4 ;
      RECT 0.000 85.412 0.140 85.552 ;
      END
    END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 84.855 0.140 84.995 ;
      LAYER metal2 ;
      RECT 0.000 84.855 0.140 84.995 ;
      LAYER metal3 ;
      RECT 0.000 84.855 0.140 84.995 ;
      LAYER metal4 ;
      RECT 0.000 84.855 0.140 84.995 ;
      END
    END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 84.297 0.140 84.437 ;
      LAYER metal2 ;
      RECT 0.000 84.297 0.140 84.437 ;
      LAYER metal3 ;
      RECT 0.000 84.297 0.140 84.437 ;
      LAYER metal4 ;
      RECT 0.000 84.297 0.140 84.437 ;
      END
    END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 83.740 0.140 83.880 ;
      LAYER metal2 ;
      RECT 0.000 83.740 0.140 83.880 ;
      LAYER metal3 ;
      RECT 0.000 83.740 0.140 83.880 ;
      LAYER metal4 ;
      RECT 0.000 83.740 0.140 83.880 ;
      END
    END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 83.183 0.140 83.323 ;
      LAYER metal2 ;
      RECT 0.000 83.183 0.140 83.323 ;
      LAYER metal3 ;
      RECT 0.000 83.183 0.140 83.323 ;
      LAYER metal4 ;
      RECT 0.000 83.183 0.140 83.323 ;
      END
    END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 82.625 0.140 82.765 ;
      LAYER metal2 ;
      RECT 0.000 82.625 0.140 82.765 ;
      LAYER metal3 ;
      RECT 0.000 82.625 0.140 82.765 ;
      LAYER metal4 ;
      RECT 0.000 82.625 0.140 82.765 ;
      END
    END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 82.068 0.140 82.208 ;
      LAYER metal2 ;
      RECT 0.000 82.068 0.140 82.208 ;
      LAYER metal3 ;
      RECT 0.000 82.068 0.140 82.208 ;
      LAYER metal4 ;
      RECT 0.000 82.068 0.140 82.208 ;
      END
    END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 81.511 0.140 81.651 ;
      LAYER metal2 ;
      RECT 0.000 81.511 0.140 81.651 ;
      LAYER metal3 ;
      RECT 0.000 81.511 0.140 81.651 ;
      LAYER metal4 ;
      RECT 0.000 81.511 0.140 81.651 ;
      END
    END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 80.954 0.140 81.094 ;
      LAYER metal2 ;
      RECT 0.000 80.954 0.140 81.094 ;
      LAYER metal3 ;
      RECT 0.000 80.954 0.140 81.094 ;
      LAYER metal4 ;
      RECT 0.000 80.954 0.140 81.094 ;
      END
    END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 80.396 0.140 80.536 ;
      LAYER metal2 ;
      RECT 0.000 80.396 0.140 80.536 ;
      LAYER metal3 ;
      RECT 0.000 80.396 0.140 80.536 ;
      LAYER metal4 ;
      RECT 0.000 80.396 0.140 80.536 ;
      END
    END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 79.839 0.140 79.979 ;
      LAYER metal2 ;
      RECT 0.000 79.839 0.140 79.979 ;
      LAYER metal3 ;
      RECT 0.000 79.839 0.140 79.979 ;
      LAYER metal4 ;
      RECT 0.000 79.839 0.140 79.979 ;
      END
    END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 79.282 0.140 79.422 ;
      LAYER metal2 ;
      RECT 0.000 79.282 0.140 79.422 ;
      LAYER metal3 ;
      RECT 0.000 79.282 0.140 79.422 ;
      LAYER metal4 ;
      RECT 0.000 79.282 0.140 79.422 ;
      END
    END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 78.724 0.140 78.864 ;
      LAYER metal2 ;
      RECT 0.000 78.724 0.140 78.864 ;
      LAYER metal3 ;
      RECT 0.000 78.724 0.140 78.864 ;
      LAYER metal4 ;
      RECT 0.000 78.724 0.140 78.864 ;
      END
    END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 78.167 0.140 78.307 ;
      LAYER metal2 ;
      RECT 0.000 78.167 0.140 78.307 ;
      LAYER metal3 ;
      RECT 0.000 78.167 0.140 78.307 ;
      LAYER metal4 ;
      RECT 0.000 78.167 0.140 78.307 ;
      END
    END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 77.610 0.140 77.750 ;
      LAYER metal2 ;
      RECT 0.000 77.610 0.140 77.750 ;
      LAYER metal3 ;
      RECT 0.000 77.610 0.140 77.750 ;
      LAYER metal4 ;
      RECT 0.000 77.610 0.140 77.750 ;
      END
    END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 77.052 0.140 77.192 ;
      LAYER metal2 ;
      RECT 0.000 77.052 0.140 77.192 ;
      LAYER metal3 ;
      RECT 0.000 77.052 0.140 77.192 ;
      LAYER metal4 ;
      RECT 0.000 77.052 0.140 77.192 ;
      END
    END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 76.495 0.140 76.635 ;
      LAYER metal2 ;
      RECT 0.000 76.495 0.140 76.635 ;
      LAYER metal3 ;
      RECT 0.000 76.495 0.140 76.635 ;
      LAYER metal4 ;
      RECT 0.000 76.495 0.140 76.635 ;
      END
    END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 75.938 0.140 76.078 ;
      LAYER metal2 ;
      RECT 0.000 75.938 0.140 76.078 ;
      LAYER metal3 ;
      RECT 0.000 75.938 0.140 76.078 ;
      LAYER metal4 ;
      RECT 0.000 75.938 0.140 76.078 ;
      END
    END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 75.381 0.140 75.521 ;
      LAYER metal2 ;
      RECT 0.000 75.381 0.140 75.521 ;
      LAYER metal3 ;
      RECT 0.000 75.381 0.140 75.521 ;
      LAYER metal4 ;
      RECT 0.000 75.381 0.140 75.521 ;
      END
    END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 74.823 0.140 74.963 ;
      LAYER metal2 ;
      RECT 0.000 74.823 0.140 74.963 ;
      LAYER metal3 ;
      RECT 0.000 74.823 0.140 74.963 ;
      LAYER metal4 ;
      RECT 0.000 74.823 0.140 74.963 ;
      END
    END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 74.266 0.140 74.406 ;
      LAYER metal2 ;
      RECT 0.000 74.266 0.140 74.406 ;
      LAYER metal3 ;
      RECT 0.000 74.266 0.140 74.406 ;
      LAYER metal4 ;
      RECT 0.000 74.266 0.140 74.406 ;
      END
    END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 73.709 0.140 73.849 ;
      LAYER metal2 ;
      RECT 0.000 73.709 0.140 73.849 ;
      LAYER metal3 ;
      RECT 0.000 73.709 0.140 73.849 ;
      LAYER metal4 ;
      RECT 0.000 73.709 0.140 73.849 ;
      END
    END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 73.151 0.140 73.291 ;
      LAYER metal2 ;
      RECT 0.000 73.151 0.140 73.291 ;
      LAYER metal3 ;
      RECT 0.000 73.151 0.140 73.291 ;
      LAYER metal4 ;
      RECT 0.000 73.151 0.140 73.291 ;
      END
    END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 72.594 0.140 72.734 ;
      LAYER metal2 ;
      RECT 0.000 72.594 0.140 72.734 ;
      LAYER metal3 ;
      RECT 0.000 72.594 0.140 72.734 ;
      LAYER metal4 ;
      RECT 0.000 72.594 0.140 72.734 ;
      END
    END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 72.037 0.140 72.177 ;
      LAYER metal2 ;
      RECT 0.000 72.037 0.140 72.177 ;
      LAYER metal3 ;
      RECT 0.000 72.037 0.140 72.177 ;
      LAYER metal4 ;
      RECT 0.000 72.037 0.140 72.177 ;
      END
    END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 71.480 0.140 71.620 ;
      LAYER metal2 ;
      RECT 0.000 71.480 0.140 71.620 ;
      LAYER metal3 ;
      RECT 0.000 71.480 0.140 71.620 ;
      LAYER metal4 ;
      RECT 0.000 71.480 0.140 71.620 ;
      END
    END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 70.922 0.140 71.062 ;
      LAYER metal2 ;
      RECT 0.000 70.922 0.140 71.062 ;
      LAYER metal3 ;
      RECT 0.000 70.922 0.140 71.062 ;
      LAYER metal4 ;
      RECT 0.000 70.922 0.140 71.062 ;
      END
    END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 70.365 0.140 70.505 ;
      LAYER metal2 ;
      RECT 0.000 70.365 0.140 70.505 ;
      LAYER metal3 ;
      RECT 0.000 70.365 0.140 70.505 ;
      LAYER metal4 ;
      RECT 0.000 70.365 0.140 70.505 ;
      END
    END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 69.808 0.140 69.948 ;
      LAYER metal2 ;
      RECT 0.000 69.808 0.140 69.948 ;
      LAYER metal3 ;
      RECT 0.000 69.808 0.140 69.948 ;
      LAYER metal4 ;
      RECT 0.000 69.808 0.140 69.948 ;
      END
    END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 69.250 0.140 69.390 ;
      LAYER metal2 ;
      RECT 0.000 69.250 0.140 69.390 ;
      LAYER metal3 ;
      RECT 0.000 69.250 0.140 69.390 ;
      LAYER metal4 ;
      RECT 0.000 69.250 0.140 69.390 ;
      END
    END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 68.693 0.140 68.833 ;
      LAYER metal2 ;
      RECT 0.000 68.693 0.140 68.833 ;
      LAYER metal3 ;
      RECT 0.000 68.693 0.140 68.833 ;
      LAYER metal4 ;
      RECT 0.000 68.693 0.140 68.833 ;
      END
    END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 68.136 0.140 68.276 ;
      LAYER metal2 ;
      RECT 0.000 68.136 0.140 68.276 ;
      LAYER metal3 ;
      RECT 0.000 68.136 0.140 68.276 ;
      LAYER metal4 ;
      RECT 0.000 68.136 0.140 68.276 ;
      END
    END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 67.578 0.140 67.718 ;
      LAYER metal2 ;
      RECT 0.000 67.578 0.140 67.718 ;
      LAYER metal3 ;
      RECT 0.000 67.578 0.140 67.718 ;
      LAYER metal4 ;
      RECT 0.000 67.578 0.140 67.718 ;
      END
    END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 67.021 0.140 67.161 ;
      LAYER metal2 ;
      RECT 0.000 67.021 0.140 67.161 ;
      LAYER metal3 ;
      RECT 0.000 67.021 0.140 67.161 ;
      LAYER metal4 ;
      RECT 0.000 67.021 0.140 67.161 ;
      END
    END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 66.464 0.140 66.604 ;
      LAYER metal2 ;
      RECT 0.000 66.464 0.140 66.604 ;
      LAYER metal3 ;
      RECT 0.000 66.464 0.140 66.604 ;
      LAYER metal4 ;
      RECT 0.000 66.464 0.140 66.604 ;
      END
    END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 65.907 0.140 66.047 ;
      LAYER metal2 ;
      RECT 0.000 65.907 0.140 66.047 ;
      LAYER metal3 ;
      RECT 0.000 65.907 0.140 66.047 ;
      LAYER metal4 ;
      RECT 0.000 65.907 0.140 66.047 ;
      END
    END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 65.349 0.140 65.489 ;
      LAYER metal2 ;
      RECT 0.000 65.349 0.140 65.489 ;
      LAYER metal3 ;
      RECT 0.000 65.349 0.140 65.489 ;
      LAYER metal4 ;
      RECT 0.000 65.349 0.140 65.489 ;
      END
    END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 64.792 0.140 64.932 ;
      LAYER metal2 ;
      RECT 0.000 64.792 0.140 64.932 ;
      LAYER metal3 ;
      RECT 0.000 64.792 0.140 64.932 ;
      LAYER metal4 ;
      RECT 0.000 64.792 0.140 64.932 ;
      END
    END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 64.235 0.140 64.375 ;
      LAYER metal2 ;
      RECT 0.000 64.235 0.140 64.375 ;
      LAYER metal3 ;
      RECT 0.000 64.235 0.140 64.375 ;
      LAYER metal4 ;
      RECT 0.000 64.235 0.140 64.375 ;
      END
    END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 63.677 0.140 63.817 ;
      LAYER metal2 ;
      RECT 0.000 63.677 0.140 63.817 ;
      LAYER metal3 ;
      RECT 0.000 63.677 0.140 63.817 ;
      LAYER metal4 ;
      RECT 0.000 63.677 0.140 63.817 ;
      END
    END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 63.120 0.140 63.260 ;
      LAYER metal2 ;
      RECT 0.000 63.120 0.140 63.260 ;
      LAYER metal3 ;
      RECT 0.000 63.120 0.140 63.260 ;
      LAYER metal4 ;
      RECT 0.000 63.120 0.140 63.260 ;
      END
    END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 62.563 0.140 62.703 ;
      LAYER metal2 ;
      RECT 0.000 62.563 0.140 62.703 ;
      LAYER metal3 ;
      RECT 0.000 62.563 0.140 62.703 ;
      LAYER metal4 ;
      RECT 0.000 62.563 0.140 62.703 ;
      END
    END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 62.005 0.140 62.145 ;
      LAYER metal2 ;
      RECT 0.000 62.005 0.140 62.145 ;
      LAYER metal3 ;
      RECT 0.000 62.005 0.140 62.145 ;
      LAYER metal4 ;
      RECT 0.000 62.005 0.140 62.145 ;
      END
    END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 61.448 0.140 61.588 ;
      LAYER metal2 ;
      RECT 0.000 61.448 0.140 61.588 ;
      LAYER metal3 ;
      RECT 0.000 61.448 0.140 61.588 ;
      LAYER metal4 ;
      RECT 0.000 61.448 0.140 61.588 ;
      END
    END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 60.891 0.140 61.031 ;
      LAYER metal2 ;
      RECT 0.000 60.891 0.140 61.031 ;
      LAYER metal3 ;
      RECT 0.000 60.891 0.140 61.031 ;
      LAYER metal4 ;
      RECT 0.000 60.891 0.140 61.031 ;
      END
    END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 60.334 0.140 60.474 ;
      LAYER metal2 ;
      RECT 0.000 60.334 0.140 60.474 ;
      LAYER metal3 ;
      RECT 0.000 60.334 0.140 60.474 ;
      LAYER metal4 ;
      RECT 0.000 60.334 0.140 60.474 ;
      END
    END rd_out[94]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 59.776 0.140 59.916 ;
      LAYER metal2 ;
      RECT 0.000 59.776 0.140 59.916 ;
      LAYER metal3 ;
      RECT 0.000 59.776 0.140 59.916 ;
      LAYER metal4 ;
      RECT 0.000 59.776 0.140 59.916 ;
      END
    END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 59.219 0.140 59.359 ;
      LAYER metal2 ;
      RECT 0.000 59.219 0.140 59.359 ;
      LAYER metal3 ;
      RECT 0.000 59.219 0.140 59.359 ;
      LAYER metal4 ;
      RECT 0.000 59.219 0.140 59.359 ;
      END
    END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 58.662 0.140 58.802 ;
      LAYER metal2 ;
      RECT 0.000 58.662 0.140 58.802 ;
      LAYER metal3 ;
      RECT 0.000 58.662 0.140 58.802 ;
      LAYER metal4 ;
      RECT 0.000 58.662 0.140 58.802 ;
      END
    END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 58.104 0.140 58.244 ;
      LAYER metal2 ;
      RECT 0.000 58.104 0.140 58.244 ;
      LAYER metal3 ;
      RECT 0.000 58.104 0.140 58.244 ;
      LAYER metal4 ;
      RECT 0.000 58.104 0.140 58.244 ;
      END
    END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 57.547 0.140 57.687 ;
      LAYER metal2 ;
      RECT 0.000 57.547 0.140 57.687 ;
      LAYER metal3 ;
      RECT 0.000 57.547 0.140 57.687 ;
      LAYER metal4 ;
      RECT 0.000 57.547 0.140 57.687 ;
      END
    END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 56.990 0.140 57.130 ;
      LAYER metal2 ;
      RECT 0.000 56.990 0.140 57.130 ;
      LAYER metal3 ;
      RECT 0.000 56.990 0.140 57.130 ;
      LAYER metal4 ;
      RECT 0.000 56.990 0.140 57.130 ;
      END
    END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 56.432 0.140 56.572 ;
      LAYER metal2 ;
      RECT 0.000 56.432 0.140 56.572 ;
      LAYER metal3 ;
      RECT 0.000 56.432 0.140 56.572 ;
      LAYER metal4 ;
      RECT 0.000 56.432 0.140 56.572 ;
      END
    END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 55.875 0.140 56.015 ;
      LAYER metal2 ;
      RECT 0.000 55.875 0.140 56.015 ;
      LAYER metal3 ;
      RECT 0.000 55.875 0.140 56.015 ;
      LAYER metal4 ;
      RECT 0.000 55.875 0.140 56.015 ;
      END
    END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 55.318 0.140 55.458 ;
      LAYER metal2 ;
      RECT 0.000 55.318 0.140 55.458 ;
      LAYER metal3 ;
      RECT 0.000 55.318 0.140 55.458 ;
      LAYER metal4 ;
      RECT 0.000 55.318 0.140 55.458 ;
      END
    END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 54.761 0.140 54.901 ;
      LAYER metal2 ;
      RECT 0.000 54.761 0.140 54.901 ;
      LAYER metal3 ;
      RECT 0.000 54.761 0.140 54.901 ;
      LAYER metal4 ;
      RECT 0.000 54.761 0.140 54.901 ;
      END
    END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 54.203 0.140 54.343 ;
      LAYER metal2 ;
      RECT 0.000 54.203 0.140 54.343 ;
      LAYER metal3 ;
      RECT 0.000 54.203 0.140 54.343 ;
      LAYER metal4 ;
      RECT 0.000 54.203 0.140 54.343 ;
      END
    END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 53.646 0.140 53.786 ;
      LAYER metal2 ;
      RECT 0.000 53.646 0.140 53.786 ;
      LAYER metal3 ;
      RECT 0.000 53.646 0.140 53.786 ;
      LAYER metal4 ;
      RECT 0.000 53.646 0.140 53.786 ;
      END
    END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 53.089 0.140 53.229 ;
      LAYER metal2 ;
      RECT 0.000 53.089 0.140 53.229 ;
      LAYER metal3 ;
      RECT 0.000 53.089 0.140 53.229 ;
      LAYER metal4 ;
      RECT 0.000 53.089 0.140 53.229 ;
      END
    END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 52.531 0.140 52.671 ;
      LAYER metal2 ;
      RECT 0.000 52.531 0.140 52.671 ;
      LAYER metal3 ;
      RECT 0.000 52.531 0.140 52.671 ;
      LAYER metal4 ;
      RECT 0.000 52.531 0.140 52.671 ;
      END
    END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 51.974 0.140 52.114 ;
      LAYER metal2 ;
      RECT 0.000 51.974 0.140 52.114 ;
      LAYER metal3 ;
      RECT 0.000 51.974 0.140 52.114 ;
      LAYER metal4 ;
      RECT 0.000 51.974 0.140 52.114 ;
      END
    END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 51.417 0.140 51.557 ;
      LAYER metal2 ;
      RECT 0.000 51.417 0.140 51.557 ;
      LAYER metal3 ;
      RECT 0.000 51.417 0.140 51.557 ;
      LAYER metal4 ;
      RECT 0.000 51.417 0.140 51.557 ;
      END
    END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 50.860 0.140 51.000 ;
      LAYER metal2 ;
      RECT 0.000 50.860 0.140 51.000 ;
      LAYER metal3 ;
      RECT 0.000 50.860 0.140 51.000 ;
      LAYER metal4 ;
      RECT 0.000 50.860 0.140 51.000 ;
      END
    END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 50.302 0.140 50.442 ;
      LAYER metal2 ;
      RECT 0.000 50.302 0.140 50.442 ;
      LAYER metal3 ;
      RECT 0.000 50.302 0.140 50.442 ;
      LAYER metal4 ;
      RECT 0.000 50.302 0.140 50.442 ;
      END
    END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 49.745 0.140 49.885 ;
      LAYER metal2 ;
      RECT 0.000 49.745 0.140 49.885 ;
      LAYER metal3 ;
      RECT 0.000 49.745 0.140 49.885 ;
      LAYER metal4 ;
      RECT 0.000 49.745 0.140 49.885 ;
      END
    END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 49.188 0.140 49.328 ;
      LAYER metal2 ;
      RECT 0.000 49.188 0.140 49.328 ;
      LAYER metal3 ;
      RECT 0.000 49.188 0.140 49.328 ;
      LAYER metal4 ;
      RECT 0.000 49.188 0.140 49.328 ;
      END
    END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 48.630 0.140 48.770 ;
      LAYER metal2 ;
      RECT 0.000 48.630 0.140 48.770 ;
      LAYER metal3 ;
      RECT 0.000 48.630 0.140 48.770 ;
      LAYER metal4 ;
      RECT 0.000 48.630 0.140 48.770 ;
      END
    END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 48.073 0.140 48.213 ;
      LAYER metal2 ;
      RECT 0.000 48.073 0.140 48.213 ;
      LAYER metal3 ;
      RECT 0.000 48.073 0.140 48.213 ;
      LAYER metal4 ;
      RECT 0.000 48.073 0.140 48.213 ;
      END
    END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 47.516 0.140 47.656 ;
      LAYER metal2 ;
      RECT 0.000 47.516 0.140 47.656 ;
      LAYER metal3 ;
      RECT 0.000 47.516 0.140 47.656 ;
      LAYER metal4 ;
      RECT 0.000 47.516 0.140 47.656 ;
      END
    END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 46.958 0.140 47.098 ;
      LAYER metal2 ;
      RECT 0.000 46.958 0.140 47.098 ;
      LAYER metal3 ;
      RECT 0.000 46.958 0.140 47.098 ;
      LAYER metal4 ;
      RECT 0.000 46.958 0.140 47.098 ;
      END
    END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 46.401 0.140 46.541 ;
      LAYER metal2 ;
      RECT 0.000 46.401 0.140 46.541 ;
      LAYER metal3 ;
      RECT 0.000 46.401 0.140 46.541 ;
      LAYER metal4 ;
      RECT 0.000 46.401 0.140 46.541 ;
      END
    END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 45.844 0.140 45.984 ;
      LAYER metal2 ;
      RECT 0.000 45.844 0.140 45.984 ;
      LAYER metal3 ;
      RECT 0.000 45.844 0.140 45.984 ;
      LAYER metal4 ;
      RECT 0.000 45.844 0.140 45.984 ;
      END
    END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 45.287 0.140 45.427 ;
      LAYER metal2 ;
      RECT 0.000 45.287 0.140 45.427 ;
      LAYER metal3 ;
      RECT 0.000 45.287 0.140 45.427 ;
      LAYER metal4 ;
      RECT 0.000 45.287 0.140 45.427 ;
      END
    END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 44.729 0.140 44.869 ;
      LAYER metal2 ;
      RECT 0.000 44.729 0.140 44.869 ;
      LAYER metal3 ;
      RECT 0.000 44.729 0.140 44.869 ;
      LAYER metal4 ;
      RECT 0.000 44.729 0.140 44.869 ;
      END
    END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 44.172 0.140 44.312 ;
      LAYER metal2 ;
      RECT 0.000 44.172 0.140 44.312 ;
      LAYER metal3 ;
      RECT 0.000 44.172 0.140 44.312 ;
      LAYER metal4 ;
      RECT 0.000 44.172 0.140 44.312 ;
      END
    END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 43.615 0.140 43.755 ;
      LAYER metal2 ;
      RECT 0.000 43.615 0.140 43.755 ;
      LAYER metal3 ;
      RECT 0.000 43.615 0.140 43.755 ;
      LAYER metal4 ;
      RECT 0.000 43.615 0.140 43.755 ;
      END
    END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 43.057 0.140 43.197 ;
      LAYER metal2 ;
      RECT 0.000 43.057 0.140 43.197 ;
      LAYER metal3 ;
      RECT 0.000 43.057 0.140 43.197 ;
      LAYER metal4 ;
      RECT 0.000 43.057 0.140 43.197 ;
      END
    END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 42.500 0.140 42.640 ;
      LAYER metal2 ;
      RECT 0.000 42.500 0.140 42.640 ;
      LAYER metal3 ;
      RECT 0.000 42.500 0.140 42.640 ;
      LAYER metal4 ;
      RECT 0.000 42.500 0.140 42.640 ;
      END
    END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 41.943 0.140 42.083 ;
      LAYER metal2 ;
      RECT 0.000 41.943 0.140 42.083 ;
      LAYER metal3 ;
      RECT 0.000 41.943 0.140 42.083 ;
      LAYER metal4 ;
      RECT 0.000 41.943 0.140 42.083 ;
      END
    END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 41.385 0.140 41.525 ;
      LAYER metal2 ;
      RECT 0.000 41.385 0.140 41.525 ;
      LAYER metal3 ;
      RECT 0.000 41.385 0.140 41.525 ;
      LAYER metal4 ;
      RECT 0.000 41.385 0.140 41.525 ;
      END
    END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 40.828 0.140 40.968 ;
      LAYER metal2 ;
      RECT 0.000 40.828 0.140 40.968 ;
      LAYER metal3 ;
      RECT 0.000 40.828 0.140 40.968 ;
      LAYER metal4 ;
      RECT 0.000 40.828 0.140 40.968 ;
      END
    END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 40.271 0.140 40.411 ;
      LAYER metal2 ;
      RECT 0.000 40.271 0.140 40.411 ;
      LAYER metal3 ;
      RECT 0.000 40.271 0.140 40.411 ;
      LAYER metal4 ;
      RECT 0.000 40.271 0.140 40.411 ;
      END
    END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 39.714 0.140 39.854 ;
      LAYER metal2 ;
      RECT 0.000 39.714 0.140 39.854 ;
      LAYER metal3 ;
      RECT 0.000 39.714 0.140 39.854 ;
      LAYER metal4 ;
      RECT 0.000 39.714 0.140 39.854 ;
      END
    END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 39.156 0.140 39.296 ;
      LAYER metal2 ;
      RECT 0.000 39.156 0.140 39.296 ;
      LAYER metal3 ;
      RECT 0.000 39.156 0.140 39.296 ;
      LAYER metal4 ;
      RECT 0.000 39.156 0.140 39.296 ;
      END
    END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 38.599 0.140 38.739 ;
      LAYER metal2 ;
      RECT 0.000 38.599 0.140 38.739 ;
      LAYER metal3 ;
      RECT 0.000 38.599 0.140 38.739 ;
      LAYER metal4 ;
      RECT 0.000 38.599 0.140 38.739 ;
      END
    END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 38.042 0.140 38.182 ;
      LAYER metal2 ;
      RECT 0.000 38.042 0.140 38.182 ;
      LAYER metal3 ;
      RECT 0.000 38.042 0.140 38.182 ;
      LAYER metal4 ;
      RECT 0.000 38.042 0.140 38.182 ;
      END
    END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 37.484 0.140 37.624 ;
      LAYER metal2 ;
      RECT 0.000 37.484 0.140 37.624 ;
      LAYER metal3 ;
      RECT 0.000 37.484 0.140 37.624 ;
      LAYER metal4 ;
      RECT 0.000 37.484 0.140 37.624 ;
      END
    END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 36.927 0.140 37.067 ;
      LAYER metal2 ;
      RECT 0.000 36.927 0.140 37.067 ;
      LAYER metal3 ;
      RECT 0.000 36.927 0.140 37.067 ;
      LAYER metal4 ;
      RECT 0.000 36.927 0.140 37.067 ;
      END
    END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 36.370 0.140 36.510 ;
      LAYER metal2 ;
      RECT 0.000 36.370 0.140 36.510 ;
      LAYER metal3 ;
      RECT 0.000 36.370 0.140 36.510 ;
      LAYER metal4 ;
      RECT 0.000 36.370 0.140 36.510 ;
      END
    END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 35.812 0.140 35.952 ;
      LAYER metal2 ;
      RECT 0.000 35.812 0.140 35.952 ;
      LAYER metal3 ;
      RECT 0.000 35.812 0.140 35.952 ;
      LAYER metal4 ;
      RECT 0.000 35.812 0.140 35.952 ;
      END
    END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 35.255 0.140 35.395 ;
      LAYER metal2 ;
      RECT 0.000 35.255 0.140 35.395 ;
      LAYER metal3 ;
      RECT 0.000 35.255 0.140 35.395 ;
      LAYER metal4 ;
      RECT 0.000 35.255 0.140 35.395 ;
      END
    END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 34.698 0.140 34.838 ;
      LAYER metal2 ;
      RECT 0.000 34.698 0.140 34.838 ;
      LAYER metal3 ;
      RECT 0.000 34.698 0.140 34.838 ;
      LAYER metal4 ;
      RECT 0.000 34.698 0.140 34.838 ;
      END
    END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 34.141 0.140 34.281 ;
      LAYER metal2 ;
      RECT 0.000 34.141 0.140 34.281 ;
      LAYER metal3 ;
      RECT 0.000 34.141 0.140 34.281 ;
      LAYER metal4 ;
      RECT 0.000 34.141 0.140 34.281 ;
      END
    END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 33.583 0.140 33.723 ;
      LAYER metal2 ;
      RECT 0.000 33.583 0.140 33.723 ;
      LAYER metal3 ;
      RECT 0.000 33.583 0.140 33.723 ;
      LAYER metal4 ;
      RECT 0.000 33.583 0.140 33.723 ;
      END
    END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 33.026 0.140 33.166 ;
      LAYER metal2 ;
      RECT 0.000 33.026 0.140 33.166 ;
      LAYER metal3 ;
      RECT 0.000 33.026 0.140 33.166 ;
      LAYER metal4 ;
      RECT 0.000 33.026 0.140 33.166 ;
      END
    END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 32.469 0.140 32.609 ;
      LAYER metal2 ;
      RECT 0.000 32.469 0.140 32.609 ;
      LAYER metal3 ;
      RECT 0.000 32.469 0.140 32.609 ;
      LAYER metal4 ;
      RECT 0.000 32.469 0.140 32.609 ;
      END
    END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 31.911 0.140 32.051 ;
      LAYER metal2 ;
      RECT 0.000 31.911 0.140 32.051 ;
      LAYER metal3 ;
      RECT 0.000 31.911 0.140 32.051 ;
      LAYER metal4 ;
      RECT 0.000 31.911 0.140 32.051 ;
      END
    END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 31.354 0.140 31.494 ;
      LAYER metal2 ;
      RECT 0.000 31.354 0.140 31.494 ;
      LAYER metal3 ;
      RECT 0.000 31.354 0.140 31.494 ;
      LAYER metal4 ;
      RECT 0.000 31.354 0.140 31.494 ;
      END
    END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 30.797 0.140 30.937 ;
      LAYER metal2 ;
      RECT 0.000 30.797 0.140 30.937 ;
      LAYER metal3 ;
      RECT 0.000 30.797 0.140 30.937 ;
      LAYER metal4 ;
      RECT 0.000 30.797 0.140 30.937 ;
      END
    END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 30.239 0.140 30.379 ;
      LAYER metal2 ;
      RECT 0.000 30.239 0.140 30.379 ;
      LAYER metal3 ;
      RECT 0.000 30.239 0.140 30.379 ;
      LAYER metal4 ;
      RECT 0.000 30.239 0.140 30.379 ;
      END
    END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 29.682 0.140 29.822 ;
      LAYER metal2 ;
      RECT 0.000 29.682 0.140 29.822 ;
      LAYER metal3 ;
      RECT 0.000 29.682 0.140 29.822 ;
      LAYER metal4 ;
      RECT 0.000 29.682 0.140 29.822 ;
      END
    END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 29.125 0.140 29.265 ;
      LAYER metal2 ;
      RECT 0.000 29.125 0.140 29.265 ;
      LAYER metal3 ;
      RECT 0.000 29.125 0.140 29.265 ;
      LAYER metal4 ;
      RECT 0.000 29.125 0.140 29.265 ;
      END
    END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 28.568 0.140 28.708 ;
      LAYER metal2 ;
      RECT 0.000 28.568 0.140 28.708 ;
      LAYER metal3 ;
      RECT 0.000 28.568 0.140 28.708 ;
      LAYER metal4 ;
      RECT 0.000 28.568 0.140 28.708 ;
      END
    END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 28.010 0.140 28.150 ;
      LAYER metal2 ;
      RECT 0.000 28.010 0.140 28.150 ;
      LAYER metal3 ;
      RECT 0.000 28.010 0.140 28.150 ;
      LAYER metal4 ;
      RECT 0.000 28.010 0.140 28.150 ;
      END
    END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 27.453 0.140 27.593 ;
      LAYER metal2 ;
      RECT 0.000 27.453 0.140 27.593 ;
      LAYER metal3 ;
      RECT 0.000 27.453 0.140 27.593 ;
      LAYER metal4 ;
      RECT 0.000 27.453 0.140 27.593 ;
      END
    END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 26.896 0.140 27.036 ;
      LAYER metal2 ;
      RECT 0.000 26.896 0.140 27.036 ;
      LAYER metal3 ;
      RECT 0.000 26.896 0.140 27.036 ;
      LAYER metal4 ;
      RECT 0.000 26.896 0.140 27.036 ;
      END
    END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 26.338 0.140 26.478 ;
      LAYER metal2 ;
      RECT 0.000 26.338 0.140 26.478 ;
      LAYER metal3 ;
      RECT 0.000 26.338 0.140 26.478 ;
      LAYER metal4 ;
      RECT 0.000 26.338 0.140 26.478 ;
      END
    END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 25.781 0.140 25.921 ;
      LAYER metal2 ;
      RECT 0.000 25.781 0.140 25.921 ;
      LAYER metal3 ;
      RECT 0.000 25.781 0.140 25.921 ;
      LAYER metal4 ;
      RECT 0.000 25.781 0.140 25.921 ;
      END
    END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 25.224 0.140 25.364 ;
      LAYER metal2 ;
      RECT 0.000 25.224 0.140 25.364 ;
      LAYER metal3 ;
      RECT 0.000 25.224 0.140 25.364 ;
      LAYER metal4 ;
      RECT 0.000 25.224 0.140 25.364 ;
      END
    END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 24.667 0.140 24.807 ;
      LAYER metal2 ;
      RECT 0.000 24.667 0.140 24.807 ;
      LAYER metal3 ;
      RECT 0.000 24.667 0.140 24.807 ;
      LAYER metal4 ;
      RECT 0.000 24.667 0.140 24.807 ;
      END
    END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 24.109 0.140 24.249 ;
      LAYER metal2 ;
      RECT 0.000 24.109 0.140 24.249 ;
      LAYER metal3 ;
      RECT 0.000 24.109 0.140 24.249 ;
      LAYER metal4 ;
      RECT 0.000 24.109 0.140 24.249 ;
      END
    END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 23.552 0.140 23.692 ;
      LAYER metal2 ;
      RECT 0.000 23.552 0.140 23.692 ;
      LAYER metal3 ;
      RECT 0.000 23.552 0.140 23.692 ;
      LAYER metal4 ;
      RECT 0.000 23.552 0.140 23.692 ;
      END
    END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 22.995 0.140 23.135 ;
      LAYER metal2 ;
      RECT 0.000 22.995 0.140 23.135 ;
      LAYER metal3 ;
      RECT 0.000 22.995 0.140 23.135 ;
      LAYER metal4 ;
      RECT 0.000 22.995 0.140 23.135 ;
      END
    END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 22.437 0.140 22.577 ;
      LAYER metal2 ;
      RECT 0.000 22.437 0.140 22.577 ;
      LAYER metal3 ;
      RECT 0.000 22.437 0.140 22.577 ;
      LAYER metal4 ;
      RECT 0.000 22.437 0.140 22.577 ;
      END
    END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 21.880 0.140 22.020 ;
      LAYER metal2 ;
      RECT 0.000 21.880 0.140 22.020 ;
      LAYER metal3 ;
      RECT 0.000 21.880 0.140 22.020 ;
      LAYER metal4 ;
      RECT 0.000 21.880 0.140 22.020 ;
      END
    END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 21.323 0.140 21.463 ;
      LAYER metal2 ;
      RECT 0.000 21.323 0.140 21.463 ;
      LAYER metal3 ;
      RECT 0.000 21.323 0.140 21.463 ;
      LAYER metal4 ;
      RECT 0.000 21.323 0.140 21.463 ;
      END
    END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 20.765 0.140 20.905 ;
      LAYER metal2 ;
      RECT 0.000 20.765 0.140 20.905 ;
      LAYER metal3 ;
      RECT 0.000 20.765 0.140 20.905 ;
      LAYER metal4 ;
      RECT 0.000 20.765 0.140 20.905 ;
      END
    END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 20.208 0.140 20.348 ;
      LAYER metal2 ;
      RECT 0.000 20.208 0.140 20.348 ;
      LAYER metal3 ;
      RECT 0.000 20.208 0.140 20.348 ;
      LAYER metal4 ;
      RECT 0.000 20.208 0.140 20.348 ;
      END
    END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 19.651 0.140 19.791 ;
      LAYER metal2 ;
      RECT 0.000 19.651 0.140 19.791 ;
      LAYER metal3 ;
      RECT 0.000 19.651 0.140 19.791 ;
      LAYER metal4 ;
      RECT 0.000 19.651 0.140 19.791 ;
      END
    END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 19.094 0.140 19.234 ;
      LAYER metal2 ;
      RECT 0.000 19.094 0.140 19.234 ;
      LAYER metal3 ;
      RECT 0.000 19.094 0.140 19.234 ;
      LAYER metal4 ;
      RECT 0.000 19.094 0.140 19.234 ;
      END
    END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 18.536 0.140 18.676 ;
      LAYER metal2 ;
      RECT 0.000 18.536 0.140 18.676 ;
      LAYER metal3 ;
      RECT 0.000 18.536 0.140 18.676 ;
      LAYER metal4 ;
      RECT 0.000 18.536 0.140 18.676 ;
      END
    END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 17.979 0.140 18.119 ;
      LAYER metal2 ;
      RECT 0.000 17.979 0.140 18.119 ;
      LAYER metal3 ;
      RECT 0.000 17.979 0.140 18.119 ;
      LAYER metal4 ;
      RECT 0.000 17.979 0.140 18.119 ;
      END
    END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 17.422 0.140 17.562 ;
      LAYER metal2 ;
      RECT 0.000 17.422 0.140 17.562 ;
      LAYER metal3 ;
      RECT 0.000 17.422 0.140 17.562 ;
      LAYER metal4 ;
      RECT 0.000 17.422 0.140 17.562 ;
      END
    END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 16.864 0.140 17.004 ;
      LAYER metal2 ;
      RECT 0.000 16.864 0.140 17.004 ;
      LAYER metal3 ;
      RECT 0.000 16.864 0.140 17.004 ;
      LAYER metal4 ;
      RECT 0.000 16.864 0.140 17.004 ;
      END
    END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 16.307 0.140 16.447 ;
      LAYER metal2 ;
      RECT 0.000 16.307 0.140 16.447 ;
      LAYER metal3 ;
      RECT 0.000 16.307 0.140 16.447 ;
      LAYER metal4 ;
      RECT 0.000 16.307 0.140 16.447 ;
      END
    END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 15.750 0.140 15.890 ;
      LAYER metal2 ;
      RECT 0.000 15.750 0.140 15.890 ;
      LAYER metal3 ;
      RECT 0.000 15.750 0.140 15.890 ;
      LAYER metal4 ;
      RECT 0.000 15.750 0.140 15.890 ;
      END
    END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 15.192 0.140 15.332 ;
      LAYER metal2 ;
      RECT 0.000 15.192 0.140 15.332 ;
      LAYER metal3 ;
      RECT 0.000 15.192 0.140 15.332 ;
      LAYER metal4 ;
      RECT 0.000 15.192 0.140 15.332 ;
      END
    END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 14.635 0.140 14.775 ;
      LAYER metal2 ;
      RECT 0.000 14.635 0.140 14.775 ;
      LAYER metal3 ;
      RECT 0.000 14.635 0.140 14.775 ;
      LAYER metal4 ;
      RECT 0.000 14.635 0.140 14.775 ;
      END
    END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 14.078 0.140 14.218 ;
      LAYER metal2 ;
      RECT 0.000 14.078 0.140 14.218 ;
      LAYER metal3 ;
      RECT 0.000 14.078 0.140 14.218 ;
      LAYER metal4 ;
      RECT 0.000 14.078 0.140 14.218 ;
      END
    END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 13.521 0.140 13.661 ;
      LAYER metal2 ;
      RECT 0.000 13.521 0.140 13.661 ;
      LAYER metal3 ;
      RECT 0.000 13.521 0.140 13.661 ;
      LAYER metal4 ;
      RECT 0.000 13.521 0.140 13.661 ;
      END
    END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 12.963 0.140 13.103 ;
      LAYER metal2 ;
      RECT 0.000 12.963 0.140 13.103 ;
      LAYER metal3 ;
      RECT 0.000 12.963 0.140 13.103 ;
      LAYER metal4 ;
      RECT 0.000 12.963 0.140 13.103 ;
      END
    END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 12.406 0.140 12.546 ;
      LAYER metal2 ;
      RECT 0.000 12.406 0.140 12.546 ;
      LAYER metal3 ;
      RECT 0.000 12.406 0.140 12.546 ;
      LAYER metal4 ;
      RECT 0.000 12.406 0.140 12.546 ;
      END
    END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 11.849 0.140 11.989 ;
      LAYER metal2 ;
      RECT 0.000 11.849 0.140 11.989 ;
      LAYER metal3 ;
      RECT 0.000 11.849 0.140 11.989 ;
      LAYER metal4 ;
      RECT 0.000 11.849 0.140 11.989 ;
      END
    END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 11.291 0.140 11.431 ;
      LAYER metal2 ;
      RECT 0.000 11.291 0.140 11.431 ;
      LAYER metal3 ;
      RECT 0.000 11.291 0.140 11.431 ;
      LAYER metal4 ;
      RECT 0.000 11.291 0.140 11.431 ;
      END
    END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 10.734 0.140 10.874 ;
      LAYER metal2 ;
      RECT 0.000 10.734 0.140 10.874 ;
      LAYER metal3 ;
      RECT 0.000 10.734 0.140 10.874 ;
      LAYER metal4 ;
      RECT 0.000 10.734 0.140 10.874 ;
      END
    END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 10.177 0.140 10.317 ;
      LAYER metal2 ;
      RECT 0.000 10.177 0.140 10.317 ;
      LAYER metal3 ;
      RECT 0.000 10.177 0.140 10.317 ;
      LAYER metal4 ;
      RECT 0.000 10.177 0.140 10.317 ;
      END
    END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 9.619 0.140 9.759 ;
      LAYER metal2 ;
      RECT 0.000 9.619 0.140 9.759 ;
      LAYER metal3 ;
      RECT 0.000 9.619 0.140 9.759 ;
      LAYER metal4 ;
      RECT 0.000 9.619 0.140 9.759 ;
      END
    END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 9.062 0.140 9.202 ;
      LAYER metal2 ;
      RECT 0.000 9.062 0.140 9.202 ;
      LAYER metal3 ;
      RECT 0.000 9.062 0.140 9.202 ;
      LAYER metal4 ;
      RECT 0.000 9.062 0.140 9.202 ;
      END
    END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 8.505 0.140 8.645 ;
      LAYER metal2 ;
      RECT 0.000 8.505 0.140 8.645 ;
      LAYER metal3 ;
      RECT 0.000 8.505 0.140 8.645 ;
      LAYER metal4 ;
      RECT 0.000 8.505 0.140 8.645 ;
      END
    END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 7.948 0.140 8.088 ;
      LAYER metal2 ;
      RECT 0.000 7.948 0.140 8.088 ;
      LAYER metal3 ;
      RECT 0.000 7.948 0.140 8.088 ;
      LAYER metal4 ;
      RECT 0.000 7.948 0.140 8.088 ;
      END
    END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 7.390 0.140 7.530 ;
      LAYER metal2 ;
      RECT 0.000 7.390 0.140 7.530 ;
      LAYER metal3 ;
      RECT 0.000 7.390 0.140 7.530 ;
      LAYER metal4 ;
      RECT 0.000 7.390 0.140 7.530 ;
      END
    END wd_in[94]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 6.833 0.140 6.973 ;
      LAYER metal2 ;
      RECT 0.000 6.833 0.140 6.973 ;
      LAYER metal3 ;
      RECT 0.000 6.833 0.140 6.973 ;
      LAYER metal4 ;
      RECT 0.000 6.833 0.140 6.973 ;
      END
    END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 6.276 0.140 6.416 ;
      LAYER metal2 ;
      RECT 0.000 6.276 0.140 6.416 ;
      LAYER metal3 ;
      RECT 0.000 6.276 0.140 6.416 ;
      LAYER metal4 ;
      RECT 0.000 6.276 0.140 6.416 ;
      END
    END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 5.718 0.140 5.858 ;
      LAYER metal2 ;
      RECT 0.000 5.718 0.140 5.858 ;
      LAYER metal3 ;
      RECT 0.000 5.718 0.140 5.858 ;
      LAYER metal4 ;
      RECT 0.000 5.718 0.140 5.858 ;
      END
    END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 5.161 0.140 5.301 ;
      LAYER metal2 ;
      RECT 0.000 5.161 0.140 5.301 ;
      LAYER metal3 ;
      RECT 0.000 5.161 0.140 5.301 ;
      LAYER metal4 ;
      RECT 0.000 5.161 0.140 5.301 ;
      END
    END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 4.604 0.140 4.744 ;
      LAYER metal2 ;
      RECT 0.000 4.604 0.140 4.744 ;
      LAYER metal3 ;
      RECT 0.000 4.604 0.140 4.744 ;
      LAYER metal4 ;
      RECT 0.000 4.604 0.140 4.744 ;
      END
    END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 4.046 0.140 4.186 ;
      LAYER metal2 ;
      RECT 0.000 4.046 0.140 4.186 ;
      LAYER metal3 ;
      RECT 0.000 4.046 0.140 4.186 ;
      LAYER metal4 ;
      RECT 0.000 4.046 0.140 4.186 ;
      END
    END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 3.489 0.140 3.629 ;
      LAYER metal2 ;
      RECT 0.000 3.489 0.140 3.629 ;
      LAYER metal3 ;
      RECT 0.000 3.489 0.140 3.629 ;
      LAYER metal4 ;
      RECT 0.000 3.489 0.140 3.629 ;
      END
    END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 2.932 0.140 3.072 ;
      LAYER metal2 ;
      RECT 0.000 2.932 0.140 3.072 ;
      LAYER metal3 ;
      RECT 0.000 2.932 0.140 3.072 ;
      LAYER metal4 ;
      RECT 0.000 2.932 0.140 3.072 ;
      END
    END addr_in[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 2.375 0.140 2.515 ;
      LAYER metal2 ;
      RECT 0.000 2.375 0.140 2.515 ;
      LAYER metal3 ;
      RECT 0.000 2.375 0.140 2.515 ;
      LAYER metal4 ;
      RECT 0.000 2.375 0.140 2.515 ;
      END
    END clk
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 1.817 0.140 1.957 ;
      LAYER metal2 ;
      RECT 0.000 1.817 0.140 1.957 ;
      LAYER metal3 ;
      RECT 0.000 1.817 0.140 1.957 ;
      LAYER metal4 ;
      RECT 0.000 1.817 0.140 1.957 ;
      END
    END ce_in
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 7.182 166.360 50.271 166.920 ;
      RECT 7.182 163.560 50.271 164.120 ;
      RECT 7.182 160.760 50.271 161.320 ;
      RECT 7.182 157.960 50.271 158.520 ;
      RECT 7.182 155.160 50.271 155.720 ;
      RECT 7.182 152.360 50.271 152.920 ;
      RECT 7.182 149.560 50.271 150.120 ;
      RECT 7.182 146.760 50.271 147.320 ;
      RECT 7.182 143.960 50.271 144.520 ;
      RECT 7.182 141.160 50.271 141.720 ;
      RECT 7.182 138.360 50.271 138.920 ;
      RECT 7.182 135.560 50.271 136.120 ;
      RECT 7.182 132.760 50.271 133.320 ;
      RECT 7.182 129.960 50.271 130.520 ;
      RECT 7.182 127.160 50.271 127.720 ;
      RECT 7.182 124.360 50.271 124.920 ;
      RECT 7.182 121.560 50.271 122.120 ;
      RECT 7.182 118.760 50.271 119.320 ;
      RECT 7.182 115.960 50.271 116.520 ;
      RECT 7.182 113.160 50.271 113.720 ;
      RECT 7.182 110.360 50.271 110.920 ;
      RECT 7.182 107.560 50.271 108.120 ;
      RECT 7.182 104.760 50.271 105.320 ;
      RECT 7.182 101.960 50.271 102.520 ;
      RECT 7.182 99.160 50.271 99.720 ;
      RECT 7.182 96.360 50.271 96.920 ;
      RECT 7.182 93.560 50.271 94.120 ;
      RECT 7.182 90.760 50.271 91.320 ;
      RECT 7.182 87.960 50.271 88.520 ;
      RECT 7.182 85.160 50.271 85.720 ;
      RECT 7.182 82.360 50.271 82.920 ;
      RECT 7.182 79.560 50.271 80.120 ;
      RECT 7.182 76.760 50.271 77.320 ;
      RECT 7.182 73.960 50.271 74.520 ;
      RECT 7.182 71.160 50.271 71.720 ;
      RECT 7.182 68.360 50.271 68.920 ;
      RECT 7.182 65.560 50.271 66.120 ;
      RECT 7.182 62.760 50.271 63.320 ;
      RECT 7.182 59.960 50.271 60.520 ;
      RECT 7.182 57.160 50.271 57.720 ;
      RECT 7.182 54.360 50.271 54.920 ;
      RECT 7.182 51.560 50.271 52.120 ;
      RECT 7.182 48.760 50.271 49.320 ;
      RECT 7.182 45.960 50.271 46.520 ;
      RECT 7.182 43.160 50.271 43.720 ;
      RECT 7.182 40.360 50.271 40.920 ;
      RECT 7.182 37.560 50.271 38.120 ;
      RECT 7.182 34.760 50.271 35.320 ;
      RECT 7.182 31.960 50.271 32.520 ;
      RECT 7.182 29.160 50.271 29.720 ;
      RECT 7.182 26.360 50.271 26.920 ;
      RECT 7.182 23.560 50.271 24.120 ;
      RECT 7.182 20.760 50.271 21.320 ;
      RECT 7.182 17.960 50.271 18.520 ;
      RECT 7.182 15.160 50.271 15.720 ;
      RECT 7.182 12.360 50.271 12.920 ;
      RECT 7.182 9.560 50.271 10.120 ;
      RECT 7.182 6.760 50.271 7.320 ;
      RECT 7.182 3.960 50.271 4.520 ;
      END
    END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 7.182 164.960 50.271 165.520 ;
      RECT 7.182 162.160 50.271 162.720 ;
      RECT 7.182 159.360 50.271 159.920 ;
      RECT 7.182 156.560 50.271 157.120 ;
      RECT 7.182 153.760 50.271 154.320 ;
      RECT 7.182 150.960 50.271 151.520 ;
      RECT 7.182 148.160 50.271 148.720 ;
      RECT 7.182 145.360 50.271 145.920 ;
      RECT 7.182 142.560 50.271 143.120 ;
      RECT 7.182 139.760 50.271 140.320 ;
      RECT 7.182 136.960 50.271 137.520 ;
      RECT 7.182 134.160 50.271 134.720 ;
      RECT 7.182 131.360 50.271 131.920 ;
      RECT 7.182 128.560 50.271 129.120 ;
      RECT 7.182 125.760 50.271 126.320 ;
      RECT 7.182 122.960 50.271 123.520 ;
      RECT 7.182 120.160 50.271 120.720 ;
      RECT 7.182 117.360 50.271 117.920 ;
      RECT 7.182 114.560 50.271 115.120 ;
      RECT 7.182 111.760 50.271 112.320 ;
      RECT 7.182 108.960 50.271 109.520 ;
      RECT 7.182 106.160 50.271 106.720 ;
      RECT 7.182 103.360 50.271 103.920 ;
      RECT 7.182 100.560 50.271 101.120 ;
      RECT 7.182 97.760 50.271 98.320 ;
      RECT 7.182 94.960 50.271 95.520 ;
      RECT 7.182 92.160 50.271 92.720 ;
      RECT 7.182 89.360 50.271 89.920 ;
      RECT 7.182 86.560 50.271 87.120 ;
      RECT 7.182 83.760 50.271 84.320 ;
      RECT 7.182 80.960 50.271 81.520 ;
      RECT 7.182 78.160 50.271 78.720 ;
      RECT 7.182 75.360 50.271 75.920 ;
      RECT 7.182 72.560 50.271 73.120 ;
      RECT 7.182 69.760 50.271 70.320 ;
      RECT 7.182 66.960 50.271 67.520 ;
      RECT 7.182 64.160 50.271 64.720 ;
      RECT 7.182 61.360 50.271 61.920 ;
      RECT 7.182 58.560 50.271 59.120 ;
      RECT 7.182 55.760 50.271 56.320 ;
      RECT 7.182 52.960 50.271 53.520 ;
      RECT 7.182 50.160 50.271 50.720 ;
      RECT 7.182 47.360 50.271 47.920 ;
      RECT 7.182 44.560 50.271 45.120 ;
      RECT 7.182 41.760 50.271 42.320 ;
      RECT 7.182 38.960 50.271 39.520 ;
      RECT 7.182 36.160 50.271 36.720 ;
      RECT 7.182 33.360 50.271 33.920 ;
      RECT 7.182 30.560 50.271 31.120 ;
      RECT 7.182 27.760 50.271 28.320 ;
      RECT 7.182 24.960 50.271 25.520 ;
      RECT 7.182 22.160 50.271 22.720 ;
      RECT 7.182 19.360 50.271 19.920 ;
      RECT 7.182 16.560 50.271 17.120 ;
      RECT 7.182 13.760 50.271 14.320 ;
      RECT 7.182 10.960 50.271 11.520 ;
      RECT 7.182 8.160 50.271 8.720 ;
      RECT 7.182 5.360 50.271 5.920 ;
      RECT 7.182 2.560 50.271 3.120 ;
      END
    END VDD
  OBS
    LAYER metal1 ;
    RECT 0.000 167.760 57.452 166.360 ;
    RECT 0.140 166.360 57.452 166.220 ;
    RECT 0.000 166.220 57.452 165.803 ;
    RECT 0.140 165.803 57.452 165.663 ;
    RECT 0.000 165.663 57.452 165.246 ;
    RECT 0.140 165.246 57.452 165.106 ;
    RECT 0.000 165.106 57.452 164.688 ;
    RECT 0.140 164.688 57.452 164.548 ;
    RECT 0.000 164.548 57.452 164.131 ;
    RECT 0.140 164.131 57.452 163.991 ;
    RECT 0.000 163.991 57.452 163.574 ;
    RECT 0.140 163.574 57.452 163.434 ;
    RECT 0.000 163.434 57.452 163.016 ;
    RECT 0.140 163.016 57.452 162.876 ;
    RECT 0.000 162.876 57.452 162.459 ;
    RECT 0.140 162.459 57.452 162.319 ;
    RECT 0.000 162.319 57.452 161.902 ;
    RECT 0.140 161.902 57.452 161.762 ;
    RECT 0.000 161.762 57.452 161.344 ;
    RECT 0.140 161.344 57.452 161.204 ;
    RECT 0.000 161.204 57.452 160.787 ;
    RECT 0.140 160.787 57.452 160.647 ;
    RECT 0.000 160.647 57.452 160.230 ;
    RECT 0.140 160.230 57.452 160.090 ;
    RECT 0.000 160.090 57.452 159.673 ;
    RECT 0.140 159.673 57.452 159.533 ;
    RECT 0.000 159.533 57.452 159.115 ;
    RECT 0.140 159.115 57.452 158.975 ;
    RECT 0.000 158.975 57.452 158.558 ;
    RECT 0.140 158.558 57.452 158.418 ;
    RECT 0.000 158.418 57.452 158.001 ;
    RECT 0.140 158.001 57.452 157.861 ;
    RECT 0.000 157.861 57.452 157.443 ;
    RECT 0.140 157.443 57.452 157.303 ;
    RECT 0.000 157.303 57.452 156.886 ;
    RECT 0.140 156.886 57.452 156.746 ;
    RECT 0.000 156.746 57.452 156.329 ;
    RECT 0.140 156.329 57.452 156.189 ;
    RECT 0.000 156.189 57.452 155.771 ;
    RECT 0.140 155.771 57.452 155.631 ;
    RECT 0.000 155.631 57.452 155.214 ;
    RECT 0.140 155.214 57.452 155.074 ;
    RECT 0.000 155.074 57.452 154.657 ;
    RECT 0.140 154.657 57.452 154.517 ;
    RECT 0.000 154.517 57.452 154.100 ;
    RECT 0.140 154.100 57.452 153.960 ;
    RECT 0.000 153.960 57.452 153.542 ;
    RECT 0.140 153.542 57.452 153.402 ;
    RECT 0.000 153.402 57.452 152.985 ;
    RECT 0.140 152.985 57.452 152.845 ;
    RECT 0.000 152.845 57.452 152.428 ;
    RECT 0.140 152.428 57.452 152.288 ;
    RECT 0.000 152.288 57.452 151.870 ;
    RECT 0.140 151.870 57.452 151.730 ;
    RECT 0.000 151.730 57.452 151.313 ;
    RECT 0.140 151.313 57.452 151.173 ;
    RECT 0.000 151.173 57.452 150.756 ;
    RECT 0.140 150.756 57.452 150.616 ;
    RECT 0.000 150.616 57.452 150.199 ;
    RECT 0.140 150.199 57.452 150.059 ;
    RECT 0.000 150.059 57.452 149.641 ;
    RECT 0.140 149.641 57.452 149.501 ;
    RECT 0.000 149.501 57.452 149.084 ;
    RECT 0.140 149.084 57.452 148.944 ;
    RECT 0.000 148.944 57.452 148.527 ;
    RECT 0.140 148.527 57.452 148.387 ;
    RECT 0.000 148.387 57.452 147.969 ;
    RECT 0.140 147.969 57.452 147.829 ;
    RECT 0.000 147.829 57.452 147.412 ;
    RECT 0.140 147.412 57.452 147.272 ;
    RECT 0.000 147.272 57.452 146.855 ;
    RECT 0.140 146.855 57.452 146.715 ;
    RECT 0.000 146.715 57.452 146.297 ;
    RECT 0.140 146.297 57.452 146.157 ;
    RECT 0.000 146.157 57.452 145.740 ;
    RECT 0.140 145.740 57.452 145.600 ;
    RECT 0.000 145.600 57.452 145.183 ;
    RECT 0.140 145.183 57.452 145.043 ;
    RECT 0.000 145.043 57.452 144.626 ;
    RECT 0.140 144.626 57.452 144.486 ;
    RECT 0.000 144.486 57.452 144.068 ;
    RECT 0.140 144.068 57.452 143.928 ;
    RECT 0.000 143.928 57.452 143.511 ;
    RECT 0.140 143.511 57.452 143.371 ;
    RECT 0.000 143.371 57.452 142.954 ;
    RECT 0.140 142.954 57.452 142.814 ;
    RECT 0.000 142.814 57.452 142.396 ;
    RECT 0.140 142.396 57.452 142.256 ;
    RECT 0.000 142.256 57.452 141.839 ;
    RECT 0.140 141.839 57.452 141.699 ;
    RECT 0.000 141.699 57.452 141.282 ;
    RECT 0.140 141.282 57.452 141.142 ;
    RECT 0.000 141.142 57.452 140.724 ;
    RECT 0.140 140.724 57.452 140.584 ;
    RECT 0.000 140.584 57.452 140.167 ;
    RECT 0.140 140.167 57.452 140.027 ;
    RECT 0.000 140.027 57.452 139.610 ;
    RECT 0.140 139.610 57.452 139.470 ;
    RECT 0.000 139.470 57.452 139.053 ;
    RECT 0.140 139.053 57.452 138.913 ;
    RECT 0.000 138.913 57.452 138.495 ;
    RECT 0.140 138.495 57.452 138.355 ;
    RECT 0.000 138.355 57.452 137.938 ;
    RECT 0.140 137.938 57.452 137.798 ;
    RECT 0.000 137.798 57.452 137.381 ;
    RECT 0.140 137.381 57.452 137.241 ;
    RECT 0.000 137.241 57.452 136.823 ;
    RECT 0.140 136.823 57.452 136.683 ;
    RECT 0.000 136.683 57.452 136.266 ;
    RECT 0.140 136.266 57.452 136.126 ;
    RECT 0.000 136.126 57.452 135.709 ;
    RECT 0.140 135.709 57.452 135.569 ;
    RECT 0.000 135.569 57.452 135.151 ;
    RECT 0.140 135.151 57.452 135.011 ;
    RECT 0.000 135.011 57.452 134.594 ;
    RECT 0.140 134.594 57.452 134.454 ;
    RECT 0.000 134.454 57.452 134.037 ;
    RECT 0.140 134.037 57.452 133.897 ;
    RECT 0.000 133.897 57.452 133.480 ;
    RECT 0.140 133.480 57.452 133.340 ;
    RECT 0.000 133.340 57.452 132.922 ;
    RECT 0.140 132.922 57.452 132.782 ;
    RECT 0.000 132.782 57.452 132.365 ;
    RECT 0.140 132.365 57.452 132.225 ;
    RECT 0.000 132.225 57.452 131.808 ;
    RECT 0.140 131.808 57.452 131.668 ;
    RECT 0.000 131.668 57.452 131.250 ;
    RECT 0.140 131.250 57.452 131.110 ;
    RECT 0.000 131.110 57.452 130.693 ;
    RECT 0.140 130.693 57.452 130.553 ;
    RECT 0.000 130.553 57.452 130.136 ;
    RECT 0.140 130.136 57.452 129.996 ;
    RECT 0.000 129.996 57.452 129.578 ;
    RECT 0.140 129.578 57.452 129.438 ;
    RECT 0.000 129.438 57.452 129.021 ;
    RECT 0.140 129.021 57.452 128.881 ;
    RECT 0.000 128.881 57.452 128.464 ;
    RECT 0.140 128.464 57.452 128.324 ;
    RECT 0.000 128.324 57.452 127.907 ;
    RECT 0.140 127.907 57.452 127.767 ;
    RECT 0.000 127.767 57.452 127.349 ;
    RECT 0.140 127.349 57.452 127.209 ;
    RECT 0.000 127.209 57.452 126.792 ;
    RECT 0.140 126.792 57.452 126.652 ;
    RECT 0.000 126.652 57.452 126.235 ;
    RECT 0.140 126.235 57.452 126.095 ;
    RECT 0.000 126.095 57.452 125.677 ;
    RECT 0.140 125.677 57.452 125.537 ;
    RECT 0.000 125.537 57.452 125.120 ;
    RECT 0.140 125.120 57.452 124.980 ;
    RECT 0.000 124.980 57.452 124.563 ;
    RECT 0.140 124.563 57.452 124.423 ;
    RECT 0.000 124.423 57.452 124.006 ;
    RECT 0.140 124.006 57.452 123.866 ;
    RECT 0.000 123.866 57.452 123.448 ;
    RECT 0.140 123.448 57.452 123.308 ;
    RECT 0.000 123.308 57.452 122.891 ;
    RECT 0.140 122.891 57.452 122.751 ;
    RECT 0.000 122.751 57.452 122.334 ;
    RECT 0.140 122.334 57.452 122.194 ;
    RECT 0.000 122.194 57.452 121.776 ;
    RECT 0.140 121.776 57.452 121.636 ;
    RECT 0.000 121.636 57.452 121.219 ;
    RECT 0.140 121.219 57.452 121.079 ;
    RECT 0.000 121.079 57.452 120.662 ;
    RECT 0.140 120.662 57.452 120.522 ;
    RECT 0.000 120.522 57.452 120.104 ;
    RECT 0.140 120.104 57.452 119.964 ;
    RECT 0.000 119.964 57.452 119.547 ;
    RECT 0.140 119.547 57.452 119.407 ;
    RECT 0.000 119.407 57.452 118.990 ;
    RECT 0.140 118.990 57.452 118.850 ;
    RECT 0.000 118.850 57.452 118.433 ;
    RECT 0.140 118.433 57.452 118.293 ;
    RECT 0.000 118.293 57.452 117.875 ;
    RECT 0.140 117.875 57.452 117.735 ;
    RECT 0.000 117.735 57.452 117.318 ;
    RECT 0.140 117.318 57.452 117.178 ;
    RECT 0.000 117.178 57.452 116.761 ;
    RECT 0.140 116.761 57.452 116.621 ;
    RECT 0.000 116.621 57.452 116.203 ;
    RECT 0.140 116.203 57.452 116.063 ;
    RECT 0.000 116.063 57.452 115.646 ;
    RECT 0.140 115.646 57.452 115.506 ;
    RECT 0.000 115.506 57.452 115.089 ;
    RECT 0.140 115.089 57.452 114.949 ;
    RECT 0.000 114.949 57.452 114.531 ;
    RECT 0.140 114.531 57.452 114.391 ;
    RECT 0.000 114.391 57.452 113.974 ;
    RECT 0.140 113.974 57.452 113.834 ;
    RECT 0.000 113.834 57.452 113.417 ;
    RECT 0.140 113.417 57.452 113.277 ;
    RECT 0.000 113.277 57.452 112.860 ;
    RECT 0.140 112.860 57.452 112.720 ;
    RECT 0.000 112.720 57.452 112.302 ;
    RECT 0.140 112.302 57.452 112.162 ;
    RECT 0.000 112.162 57.452 111.745 ;
    RECT 0.140 111.745 57.452 111.605 ;
    RECT 0.000 111.605 57.452 111.188 ;
    RECT 0.140 111.188 57.452 111.048 ;
    RECT 0.000 111.048 57.452 110.630 ;
    RECT 0.140 110.630 57.452 110.490 ;
    RECT 0.000 110.490 57.452 110.073 ;
    RECT 0.140 110.073 57.452 109.933 ;
    RECT 0.000 109.933 57.452 109.516 ;
    RECT 0.140 109.516 57.452 109.376 ;
    RECT 0.000 109.376 57.452 108.958 ;
    RECT 0.140 108.958 57.452 108.818 ;
    RECT 0.000 108.818 57.452 108.401 ;
    RECT 0.140 108.401 57.452 108.261 ;
    RECT 0.000 108.261 57.452 107.844 ;
    RECT 0.140 107.844 57.452 107.704 ;
    RECT 0.000 107.704 57.452 107.287 ;
    RECT 0.140 107.287 57.452 107.147 ;
    RECT 0.000 107.147 57.452 106.729 ;
    RECT 0.140 106.729 57.452 106.589 ;
    RECT 0.000 106.589 57.452 106.172 ;
    RECT 0.140 106.172 57.452 106.032 ;
    RECT 0.000 106.032 57.452 105.615 ;
    RECT 0.140 105.615 57.452 105.475 ;
    RECT 0.000 105.475 57.452 105.057 ;
    RECT 0.140 105.057 57.452 104.917 ;
    RECT 0.000 104.917 57.452 104.500 ;
    RECT 0.140 104.500 57.452 104.360 ;
    RECT 0.000 104.360 57.452 103.943 ;
    RECT 0.140 103.943 57.452 103.803 ;
    RECT 0.000 103.803 57.452 103.385 ;
    RECT 0.140 103.385 57.452 103.245 ;
    RECT 0.000 103.245 57.452 102.828 ;
    RECT 0.140 102.828 57.452 102.688 ;
    RECT 0.000 102.688 57.452 102.271 ;
    RECT 0.140 102.271 57.452 102.131 ;
    RECT 0.000 102.131 57.452 101.714 ;
    RECT 0.140 101.714 57.452 101.574 ;
    RECT 0.000 101.574 57.452 101.156 ;
    RECT 0.140 101.156 57.452 101.016 ;
    RECT 0.000 101.016 57.452 100.599 ;
    RECT 0.140 100.599 57.452 100.459 ;
    RECT 0.000 100.459 57.452 100.042 ;
    RECT 0.140 100.042 57.452 99.902 ;
    RECT 0.000 99.902 57.452 99.484 ;
    RECT 0.140 99.484 57.452 99.344 ;
    RECT 0.000 99.344 57.452 98.927 ;
    RECT 0.140 98.927 57.452 98.787 ;
    RECT 0.000 98.787 57.452 98.370 ;
    RECT 0.140 98.370 57.452 98.230 ;
    RECT 0.000 98.230 57.452 97.813 ;
    RECT 0.140 97.813 57.452 97.673 ;
    RECT 0.000 97.673 57.452 97.255 ;
    RECT 0.140 97.255 57.452 97.115 ;
    RECT 0.000 97.115 57.452 96.698 ;
    RECT 0.140 96.698 57.452 96.558 ;
    RECT 0.000 96.558 57.452 96.141 ;
    RECT 0.140 96.141 57.452 96.001 ;
    RECT 0.000 96.001 57.452 95.583 ;
    RECT 0.140 95.583 57.452 95.443 ;
    RECT 0.000 95.443 57.452 95.026 ;
    RECT 0.140 95.026 57.452 94.886 ;
    RECT 0.000 94.886 57.452 94.469 ;
    RECT 0.140 94.469 57.452 94.329 ;
    RECT 0.000 94.329 57.452 93.911 ;
    RECT 0.140 93.911 57.452 93.771 ;
    RECT 0.000 93.771 57.452 93.354 ;
    RECT 0.140 93.354 57.452 93.214 ;
    RECT 0.000 93.214 57.452 92.797 ;
    RECT 0.140 92.797 57.452 92.657 ;
    RECT 0.000 92.657 57.452 92.240 ;
    RECT 0.140 92.240 57.452 92.100 ;
    RECT 0.000 92.100 57.452 91.682 ;
    RECT 0.140 91.682 57.452 91.542 ;
    RECT 0.000 91.542 57.452 91.125 ;
    RECT 0.140 91.125 57.452 90.985 ;
    RECT 0.000 90.985 57.452 90.568 ;
    RECT 0.140 90.568 57.452 90.428 ;
    RECT 0.000 90.428 57.452 90.010 ;
    RECT 0.140 90.010 57.452 89.870 ;
    RECT 0.000 89.870 57.452 89.453 ;
    RECT 0.140 89.453 57.452 89.313 ;
    RECT 0.000 89.313 57.452 88.896 ;
    RECT 0.140 88.896 57.452 88.756 ;
    RECT 0.000 88.756 57.452 88.338 ;
    RECT 0.140 88.338 57.452 88.198 ;
    RECT 0.000 88.198 57.452 87.781 ;
    RECT 0.140 87.781 57.452 87.641 ;
    RECT 0.000 87.641 57.452 87.224 ;
    RECT 0.140 87.224 57.452 87.084 ;
    RECT 0.000 87.084 57.452 86.667 ;
    RECT 0.140 86.667 57.452 86.527 ;
    RECT 0.000 86.527 57.452 86.109 ;
    RECT 0.140 86.109 57.452 85.969 ;
    RECT 0.000 85.969 57.452 85.552 ;
    RECT 0.140 85.552 57.452 85.412 ;
    RECT 0.000 85.412 57.452 84.995 ;
    RECT 0.140 84.995 57.452 84.855 ;
    RECT 0.000 84.855 57.452 84.437 ;
    RECT 0.140 84.437 57.452 84.297 ;
    RECT 0.000 84.297 57.452 83.880 ;
    RECT 0.140 83.880 57.452 83.740 ;
    RECT 0.000 83.740 57.452 83.323 ;
    RECT 0.140 83.323 57.452 83.183 ;
    RECT 0.000 83.183 57.452 82.765 ;
    RECT 0.140 82.765 57.452 82.625 ;
    RECT 0.000 82.625 57.452 82.208 ;
    RECT 0.140 82.208 57.452 82.068 ;
    RECT 0.000 82.068 57.452 81.651 ;
    RECT 0.140 81.651 57.452 81.511 ;
    RECT 0.000 81.511 57.452 81.094 ;
    RECT 0.140 81.094 57.452 80.954 ;
    RECT 0.000 80.954 57.452 80.536 ;
    RECT 0.140 80.536 57.452 80.396 ;
    RECT 0.000 80.396 57.452 79.979 ;
    RECT 0.140 79.979 57.452 79.839 ;
    RECT 0.000 79.839 57.452 79.422 ;
    RECT 0.140 79.422 57.452 79.282 ;
    RECT 0.000 79.282 57.452 78.864 ;
    RECT 0.140 78.864 57.452 78.724 ;
    RECT 0.000 78.724 57.452 78.307 ;
    RECT 0.140 78.307 57.452 78.167 ;
    RECT 0.000 78.167 57.452 77.750 ;
    RECT 0.140 77.750 57.452 77.610 ;
    RECT 0.000 77.610 57.452 77.192 ;
    RECT 0.140 77.192 57.452 77.052 ;
    RECT 0.000 77.052 57.452 76.635 ;
    RECT 0.140 76.635 57.452 76.495 ;
    RECT 0.000 76.495 57.452 76.078 ;
    RECT 0.140 76.078 57.452 75.938 ;
    RECT 0.000 75.938 57.452 75.521 ;
    RECT 0.140 75.521 57.452 75.381 ;
    RECT 0.000 75.381 57.452 74.963 ;
    RECT 0.140 74.963 57.452 74.823 ;
    RECT 0.000 74.823 57.452 74.406 ;
    RECT 0.140 74.406 57.452 74.266 ;
    RECT 0.000 74.266 57.452 73.849 ;
    RECT 0.140 73.849 57.452 73.709 ;
    RECT 0.000 73.709 57.452 73.291 ;
    RECT 0.140 73.291 57.452 73.151 ;
    RECT 0.000 73.151 57.452 72.734 ;
    RECT 0.140 72.734 57.452 72.594 ;
    RECT 0.000 72.594 57.452 72.177 ;
    RECT 0.140 72.177 57.452 72.037 ;
    RECT 0.000 72.037 57.452 71.620 ;
    RECT 0.140 71.620 57.452 71.480 ;
    RECT 0.000 71.480 57.452 71.062 ;
    RECT 0.140 71.062 57.452 70.922 ;
    RECT 0.000 70.922 57.452 70.505 ;
    RECT 0.140 70.505 57.452 70.365 ;
    RECT 0.000 70.365 57.452 69.948 ;
    RECT 0.140 69.948 57.452 69.808 ;
    RECT 0.000 69.808 57.452 69.390 ;
    RECT 0.140 69.390 57.452 69.250 ;
    RECT 0.000 69.250 57.452 68.833 ;
    RECT 0.140 68.833 57.452 68.693 ;
    RECT 0.000 68.693 57.452 68.276 ;
    RECT 0.140 68.276 57.452 68.136 ;
    RECT 0.000 68.136 57.452 67.718 ;
    RECT 0.140 67.718 57.452 67.578 ;
    RECT 0.000 67.578 57.452 67.161 ;
    RECT 0.140 67.161 57.452 67.021 ;
    RECT 0.000 67.021 57.452 66.604 ;
    RECT 0.140 66.604 57.452 66.464 ;
    RECT 0.000 66.464 57.452 66.047 ;
    RECT 0.140 66.047 57.452 65.907 ;
    RECT 0.000 65.907 57.452 65.489 ;
    RECT 0.140 65.489 57.452 65.349 ;
    RECT 0.000 65.349 57.452 64.932 ;
    RECT 0.140 64.932 57.452 64.792 ;
    RECT 0.000 64.792 57.452 64.375 ;
    RECT 0.140 64.375 57.452 64.235 ;
    RECT 0.000 64.235 57.452 63.817 ;
    RECT 0.140 63.817 57.452 63.677 ;
    RECT 0.000 63.677 57.452 63.260 ;
    RECT 0.140 63.260 57.452 63.120 ;
    RECT 0.000 63.120 57.452 62.703 ;
    RECT 0.140 62.703 57.452 62.563 ;
    RECT 0.000 62.563 57.452 62.145 ;
    RECT 0.140 62.145 57.452 62.005 ;
    RECT 0.000 62.005 57.452 61.588 ;
    RECT 0.140 61.588 57.452 61.448 ;
    RECT 0.000 61.448 57.452 61.031 ;
    RECT 0.140 61.031 57.452 60.891 ;
    RECT 0.000 60.891 57.452 60.474 ;
    RECT 0.140 60.474 57.452 60.334 ;
    RECT 0.000 60.334 57.452 59.916 ;
    RECT 0.140 59.916 57.452 59.776 ;
    RECT 0.000 59.776 57.452 59.359 ;
    RECT 0.140 59.359 57.452 59.219 ;
    RECT 0.000 59.219 57.452 58.802 ;
    RECT 0.140 58.802 57.452 58.662 ;
    RECT 0.000 58.662 57.452 58.244 ;
    RECT 0.140 58.244 57.452 58.104 ;
    RECT 0.000 58.104 57.452 57.687 ;
    RECT 0.140 57.687 57.452 57.547 ;
    RECT 0.000 57.547 57.452 57.130 ;
    RECT 0.140 57.130 57.452 56.990 ;
    RECT 0.000 56.990 57.452 56.572 ;
    RECT 0.140 56.572 57.452 56.432 ;
    RECT 0.000 56.432 57.452 56.015 ;
    RECT 0.140 56.015 57.452 55.875 ;
    RECT 0.000 55.875 57.452 55.458 ;
    RECT 0.140 55.458 57.452 55.318 ;
    RECT 0.000 55.318 57.452 54.901 ;
    RECT 0.140 54.901 57.452 54.761 ;
    RECT 0.000 54.761 57.452 54.343 ;
    RECT 0.140 54.343 57.452 54.203 ;
    RECT 0.000 54.203 57.452 53.786 ;
    RECT 0.140 53.786 57.452 53.646 ;
    RECT 0.000 53.646 57.452 53.229 ;
    RECT 0.140 53.229 57.452 53.089 ;
    RECT 0.000 53.089 57.452 52.671 ;
    RECT 0.140 52.671 57.452 52.531 ;
    RECT 0.000 52.531 57.452 52.114 ;
    RECT 0.140 52.114 57.452 51.974 ;
    RECT 0.000 51.974 57.452 51.557 ;
    RECT 0.140 51.557 57.452 51.417 ;
    RECT 0.000 51.417 57.452 51.000 ;
    RECT 0.140 51.000 57.452 50.860 ;
    RECT 0.000 50.860 57.452 50.442 ;
    RECT 0.140 50.442 57.452 50.302 ;
    RECT 0.000 50.302 57.452 49.885 ;
    RECT 0.140 49.885 57.452 49.745 ;
    RECT 0.000 49.745 57.452 49.328 ;
    RECT 0.140 49.328 57.452 49.188 ;
    RECT 0.000 49.188 57.452 48.770 ;
    RECT 0.140 48.770 57.452 48.630 ;
    RECT 0.000 48.630 57.452 48.213 ;
    RECT 0.140 48.213 57.452 48.073 ;
    RECT 0.000 48.073 57.452 47.656 ;
    RECT 0.140 47.656 57.452 47.516 ;
    RECT 0.000 47.516 57.452 47.098 ;
    RECT 0.140 47.098 57.452 46.958 ;
    RECT 0.000 46.958 57.452 46.541 ;
    RECT 0.140 46.541 57.452 46.401 ;
    RECT 0.000 46.401 57.452 45.984 ;
    RECT 0.140 45.984 57.452 45.844 ;
    RECT 0.000 45.844 57.452 45.427 ;
    RECT 0.140 45.427 57.452 45.287 ;
    RECT 0.000 45.287 57.452 44.869 ;
    RECT 0.140 44.869 57.452 44.729 ;
    RECT 0.000 44.729 57.452 44.312 ;
    RECT 0.140 44.312 57.452 44.172 ;
    RECT 0.000 44.172 57.452 43.755 ;
    RECT 0.140 43.755 57.452 43.615 ;
    RECT 0.000 43.615 57.452 43.197 ;
    RECT 0.140 43.197 57.452 43.057 ;
    RECT 0.000 43.057 57.452 42.640 ;
    RECT 0.140 42.640 57.452 42.500 ;
    RECT 0.000 42.500 57.452 42.083 ;
    RECT 0.140 42.083 57.452 41.943 ;
    RECT 0.000 41.943 57.452 41.525 ;
    RECT 0.140 41.525 57.452 41.385 ;
    RECT 0.000 41.385 57.452 40.968 ;
    RECT 0.140 40.968 57.452 40.828 ;
    RECT 0.000 40.828 57.452 40.411 ;
    RECT 0.140 40.411 57.452 40.271 ;
    RECT 0.000 40.271 57.452 39.854 ;
    RECT 0.140 39.854 57.452 39.714 ;
    RECT 0.000 39.714 57.452 39.296 ;
    RECT 0.140 39.296 57.452 39.156 ;
    RECT 0.000 39.156 57.452 38.739 ;
    RECT 0.140 38.739 57.452 38.599 ;
    RECT 0.000 38.599 57.452 38.182 ;
    RECT 0.140 38.182 57.452 38.042 ;
    RECT 0.000 38.042 57.452 37.624 ;
    RECT 0.140 37.624 57.452 37.484 ;
    RECT 0.000 37.484 57.452 37.067 ;
    RECT 0.140 37.067 57.452 36.927 ;
    RECT 0.000 36.927 57.452 36.510 ;
    RECT 0.140 36.510 57.452 36.370 ;
    RECT 0.000 36.370 57.452 35.952 ;
    RECT 0.140 35.952 57.452 35.812 ;
    RECT 0.000 35.812 57.452 35.395 ;
    RECT 0.140 35.395 57.452 35.255 ;
    RECT 0.000 35.255 57.452 34.838 ;
    RECT 0.140 34.838 57.452 34.698 ;
    RECT 0.000 34.698 57.452 34.281 ;
    RECT 0.140 34.281 57.452 34.141 ;
    RECT 0.000 34.141 57.452 33.723 ;
    RECT 0.140 33.723 57.452 33.583 ;
    RECT 0.000 33.583 57.452 33.166 ;
    RECT 0.140 33.166 57.452 33.026 ;
    RECT 0.000 33.026 57.452 32.609 ;
    RECT 0.140 32.609 57.452 32.469 ;
    RECT 0.000 32.469 57.452 32.051 ;
    RECT 0.140 32.051 57.452 31.911 ;
    RECT 0.000 31.911 57.452 31.494 ;
    RECT 0.140 31.494 57.452 31.354 ;
    RECT 0.000 31.354 57.452 30.937 ;
    RECT 0.140 30.937 57.452 30.797 ;
    RECT 0.000 30.797 57.452 30.379 ;
    RECT 0.140 30.379 57.452 30.239 ;
    RECT 0.000 30.239 57.452 29.822 ;
    RECT 0.140 29.822 57.452 29.682 ;
    RECT 0.000 29.682 57.452 29.265 ;
    RECT 0.140 29.265 57.452 29.125 ;
    RECT 0.000 29.125 57.452 28.708 ;
    RECT 0.140 28.708 57.452 28.568 ;
    RECT 0.000 28.568 57.452 28.150 ;
    RECT 0.140 28.150 57.452 28.010 ;
    RECT 0.000 28.010 57.452 27.593 ;
    RECT 0.140 27.593 57.452 27.453 ;
    RECT 0.000 27.453 57.452 27.036 ;
    RECT 0.140 27.036 57.452 26.896 ;
    RECT 0.000 26.896 57.452 26.478 ;
    RECT 0.140 26.478 57.452 26.338 ;
    RECT 0.000 26.338 57.452 25.921 ;
    RECT 0.140 25.921 57.452 25.781 ;
    RECT 0.000 25.781 57.452 25.364 ;
    RECT 0.140 25.364 57.452 25.224 ;
    RECT 0.000 25.224 57.452 24.807 ;
    RECT 0.140 24.807 57.452 24.667 ;
    RECT 0.000 24.667 57.452 24.249 ;
    RECT 0.140 24.249 57.452 24.109 ;
    RECT 0.000 24.109 57.452 23.692 ;
    RECT 0.140 23.692 57.452 23.552 ;
    RECT 0.000 23.552 57.452 23.135 ;
    RECT 0.140 23.135 57.452 22.995 ;
    RECT 0.000 22.995 57.452 22.577 ;
    RECT 0.140 22.577 57.452 22.437 ;
    RECT 0.000 22.437 57.452 22.020 ;
    RECT 0.140 22.020 57.452 21.880 ;
    RECT 0.000 21.880 57.452 21.463 ;
    RECT 0.140 21.463 57.452 21.323 ;
    RECT 0.000 21.323 57.452 20.905 ;
    RECT 0.140 20.905 57.452 20.765 ;
    RECT 0.000 20.765 57.452 20.348 ;
    RECT 0.140 20.348 57.452 20.208 ;
    RECT 0.000 20.208 57.452 19.791 ;
    RECT 0.140 19.791 57.452 19.651 ;
    RECT 0.000 19.651 57.452 19.234 ;
    RECT 0.140 19.234 57.452 19.094 ;
    RECT 0.000 19.094 57.452 18.676 ;
    RECT 0.140 18.676 57.452 18.536 ;
    RECT 0.000 18.536 57.452 18.119 ;
    RECT 0.140 18.119 57.452 17.979 ;
    RECT 0.000 17.979 57.452 17.562 ;
    RECT 0.140 17.562 57.452 17.422 ;
    RECT 0.000 17.422 57.452 17.004 ;
    RECT 0.140 17.004 57.452 16.864 ;
    RECT 0.000 16.864 57.452 16.447 ;
    RECT 0.140 16.447 57.452 16.307 ;
    RECT 0.000 16.307 57.452 15.890 ;
    RECT 0.140 15.890 57.452 15.750 ;
    RECT 0.000 15.750 57.452 15.332 ;
    RECT 0.140 15.332 57.452 15.192 ;
    RECT 0.000 15.192 57.452 14.775 ;
    RECT 0.140 14.775 57.452 14.635 ;
    RECT 0.000 14.635 57.452 14.218 ;
    RECT 0.140 14.218 57.452 14.078 ;
    RECT 0.000 14.078 57.452 13.661 ;
    RECT 0.140 13.661 57.452 13.521 ;
    RECT 0.000 13.521 57.452 13.103 ;
    RECT 0.140 13.103 57.452 12.963 ;
    RECT 0.000 12.963 57.452 12.546 ;
    RECT 0.140 12.546 57.452 12.406 ;
    RECT 0.000 12.406 57.452 11.989 ;
    RECT 0.140 11.989 57.452 11.849 ;
    RECT 0.000 11.849 57.452 11.431 ;
    RECT 0.140 11.431 57.452 11.291 ;
    RECT 0.000 11.291 57.452 10.874 ;
    RECT 0.140 10.874 57.452 10.734 ;
    RECT 0.000 10.734 57.452 10.317 ;
    RECT 0.140 10.317 57.452 10.177 ;
    RECT 0.000 10.177 57.452 9.759 ;
    RECT 0.140 9.759 57.452 9.619 ;
    RECT 0.000 9.619 57.452 9.202 ;
    RECT 0.140 9.202 57.452 9.062 ;
    RECT 0.000 9.062 57.452 8.645 ;
    RECT 0.140 8.645 57.452 8.505 ;
    RECT 0.000 8.505 57.452 8.088 ;
    RECT 0.140 8.088 57.452 7.948 ;
    RECT 0.000 7.948 57.452 7.530 ;
    RECT 0.140 7.530 57.452 7.390 ;
    RECT 0.000 7.390 57.452 6.973 ;
    RECT 0.140 6.973 57.452 6.833 ;
    RECT 0.000 6.833 57.452 6.416 ;
    RECT 0.140 6.416 57.452 6.276 ;
    RECT 0.000 6.276 57.452 5.858 ;
    RECT 0.140 5.858 57.452 5.718 ;
    RECT 0.000 5.718 57.452 5.301 ;
    RECT 0.140 5.301 57.452 5.161 ;
    RECT 0.000 5.161 57.452 4.744 ;
    RECT 0.140 4.744 57.452 4.604 ;
    RECT 0.000 4.604 57.452 4.186 ;
    RECT 0.140 4.186 57.452 4.046 ;
    RECT 0.000 4.046 57.452 3.629 ;
    RECT 0.140 3.629 57.452 3.489 ;
    RECT 0.000 3.489 57.452 3.072 ;
    RECT 0.140 3.072 57.452 2.932 ;
    RECT 0.000 2.932 57.452 2.515 ;
    RECT 0.140 2.515 57.452 2.375 ;
    RECT 0.000 2.375 57.452 1.957 ;
    RECT 0.140 1.957 57.452 1.817 ;
    RECT 0.000 1.817 57.452 1.400 ;
    RECT 0.000 1.400 57.452 0.000 ;
    LAYER metal2 ;
    RECT 0.000 167.760 57.452 166.360 ;
    RECT 0.140 166.360 57.452 166.220 ;
    RECT 0.000 166.220 57.452 165.803 ;
    RECT 0.140 165.803 57.452 165.663 ;
    RECT 0.000 165.663 57.452 165.246 ;
    RECT 0.140 165.246 57.452 165.106 ;
    RECT 0.000 165.106 57.452 164.688 ;
    RECT 0.140 164.688 57.452 164.548 ;
    RECT 0.000 164.548 57.452 164.131 ;
    RECT 0.140 164.131 57.452 163.991 ;
    RECT 0.000 163.991 57.452 163.574 ;
    RECT 0.140 163.574 57.452 163.434 ;
    RECT 0.000 163.434 57.452 163.016 ;
    RECT 0.140 163.016 57.452 162.876 ;
    RECT 0.000 162.876 57.452 162.459 ;
    RECT 0.140 162.459 57.452 162.319 ;
    RECT 0.000 162.319 57.452 161.902 ;
    RECT 0.140 161.902 57.452 161.762 ;
    RECT 0.000 161.762 57.452 161.344 ;
    RECT 0.140 161.344 57.452 161.204 ;
    RECT 0.000 161.204 57.452 160.787 ;
    RECT 0.140 160.787 57.452 160.647 ;
    RECT 0.000 160.647 57.452 160.230 ;
    RECT 0.140 160.230 57.452 160.090 ;
    RECT 0.000 160.090 57.452 159.673 ;
    RECT 0.140 159.673 57.452 159.533 ;
    RECT 0.000 159.533 57.452 159.115 ;
    RECT 0.140 159.115 57.452 158.975 ;
    RECT 0.000 158.975 57.452 158.558 ;
    RECT 0.140 158.558 57.452 158.418 ;
    RECT 0.000 158.418 57.452 158.001 ;
    RECT 0.140 158.001 57.452 157.861 ;
    RECT 0.000 157.861 57.452 157.443 ;
    RECT 0.140 157.443 57.452 157.303 ;
    RECT 0.000 157.303 57.452 156.886 ;
    RECT 0.140 156.886 57.452 156.746 ;
    RECT 0.000 156.746 57.452 156.329 ;
    RECT 0.140 156.329 57.452 156.189 ;
    RECT 0.000 156.189 57.452 155.771 ;
    RECT 0.140 155.771 57.452 155.631 ;
    RECT 0.000 155.631 57.452 155.214 ;
    RECT 0.140 155.214 57.452 155.074 ;
    RECT 0.000 155.074 57.452 154.657 ;
    RECT 0.140 154.657 57.452 154.517 ;
    RECT 0.000 154.517 57.452 154.100 ;
    RECT 0.140 154.100 57.452 153.960 ;
    RECT 0.000 153.960 57.452 153.542 ;
    RECT 0.140 153.542 57.452 153.402 ;
    RECT 0.000 153.402 57.452 152.985 ;
    RECT 0.140 152.985 57.452 152.845 ;
    RECT 0.000 152.845 57.452 152.428 ;
    RECT 0.140 152.428 57.452 152.288 ;
    RECT 0.000 152.288 57.452 151.870 ;
    RECT 0.140 151.870 57.452 151.730 ;
    RECT 0.000 151.730 57.452 151.313 ;
    RECT 0.140 151.313 57.452 151.173 ;
    RECT 0.000 151.173 57.452 150.756 ;
    RECT 0.140 150.756 57.452 150.616 ;
    RECT 0.000 150.616 57.452 150.199 ;
    RECT 0.140 150.199 57.452 150.059 ;
    RECT 0.000 150.059 57.452 149.641 ;
    RECT 0.140 149.641 57.452 149.501 ;
    RECT 0.000 149.501 57.452 149.084 ;
    RECT 0.140 149.084 57.452 148.944 ;
    RECT 0.000 148.944 57.452 148.527 ;
    RECT 0.140 148.527 57.452 148.387 ;
    RECT 0.000 148.387 57.452 147.969 ;
    RECT 0.140 147.969 57.452 147.829 ;
    RECT 0.000 147.829 57.452 147.412 ;
    RECT 0.140 147.412 57.452 147.272 ;
    RECT 0.000 147.272 57.452 146.855 ;
    RECT 0.140 146.855 57.452 146.715 ;
    RECT 0.000 146.715 57.452 146.297 ;
    RECT 0.140 146.297 57.452 146.157 ;
    RECT 0.000 146.157 57.452 145.740 ;
    RECT 0.140 145.740 57.452 145.600 ;
    RECT 0.000 145.600 57.452 145.183 ;
    RECT 0.140 145.183 57.452 145.043 ;
    RECT 0.000 145.043 57.452 144.626 ;
    RECT 0.140 144.626 57.452 144.486 ;
    RECT 0.000 144.486 57.452 144.068 ;
    RECT 0.140 144.068 57.452 143.928 ;
    RECT 0.000 143.928 57.452 143.511 ;
    RECT 0.140 143.511 57.452 143.371 ;
    RECT 0.000 143.371 57.452 142.954 ;
    RECT 0.140 142.954 57.452 142.814 ;
    RECT 0.000 142.814 57.452 142.396 ;
    RECT 0.140 142.396 57.452 142.256 ;
    RECT 0.000 142.256 57.452 141.839 ;
    RECT 0.140 141.839 57.452 141.699 ;
    RECT 0.000 141.699 57.452 141.282 ;
    RECT 0.140 141.282 57.452 141.142 ;
    RECT 0.000 141.142 57.452 140.724 ;
    RECT 0.140 140.724 57.452 140.584 ;
    RECT 0.000 140.584 57.452 140.167 ;
    RECT 0.140 140.167 57.452 140.027 ;
    RECT 0.000 140.027 57.452 139.610 ;
    RECT 0.140 139.610 57.452 139.470 ;
    RECT 0.000 139.470 57.452 139.053 ;
    RECT 0.140 139.053 57.452 138.913 ;
    RECT 0.000 138.913 57.452 138.495 ;
    RECT 0.140 138.495 57.452 138.355 ;
    RECT 0.000 138.355 57.452 137.938 ;
    RECT 0.140 137.938 57.452 137.798 ;
    RECT 0.000 137.798 57.452 137.381 ;
    RECT 0.140 137.381 57.452 137.241 ;
    RECT 0.000 137.241 57.452 136.823 ;
    RECT 0.140 136.823 57.452 136.683 ;
    RECT 0.000 136.683 57.452 136.266 ;
    RECT 0.140 136.266 57.452 136.126 ;
    RECT 0.000 136.126 57.452 135.709 ;
    RECT 0.140 135.709 57.452 135.569 ;
    RECT 0.000 135.569 57.452 135.151 ;
    RECT 0.140 135.151 57.452 135.011 ;
    RECT 0.000 135.011 57.452 134.594 ;
    RECT 0.140 134.594 57.452 134.454 ;
    RECT 0.000 134.454 57.452 134.037 ;
    RECT 0.140 134.037 57.452 133.897 ;
    RECT 0.000 133.897 57.452 133.480 ;
    RECT 0.140 133.480 57.452 133.340 ;
    RECT 0.000 133.340 57.452 132.922 ;
    RECT 0.140 132.922 57.452 132.782 ;
    RECT 0.000 132.782 57.452 132.365 ;
    RECT 0.140 132.365 57.452 132.225 ;
    RECT 0.000 132.225 57.452 131.808 ;
    RECT 0.140 131.808 57.452 131.668 ;
    RECT 0.000 131.668 57.452 131.250 ;
    RECT 0.140 131.250 57.452 131.110 ;
    RECT 0.000 131.110 57.452 130.693 ;
    RECT 0.140 130.693 57.452 130.553 ;
    RECT 0.000 130.553 57.452 130.136 ;
    RECT 0.140 130.136 57.452 129.996 ;
    RECT 0.000 129.996 57.452 129.578 ;
    RECT 0.140 129.578 57.452 129.438 ;
    RECT 0.000 129.438 57.452 129.021 ;
    RECT 0.140 129.021 57.452 128.881 ;
    RECT 0.000 128.881 57.452 128.464 ;
    RECT 0.140 128.464 57.452 128.324 ;
    RECT 0.000 128.324 57.452 127.907 ;
    RECT 0.140 127.907 57.452 127.767 ;
    RECT 0.000 127.767 57.452 127.349 ;
    RECT 0.140 127.349 57.452 127.209 ;
    RECT 0.000 127.209 57.452 126.792 ;
    RECT 0.140 126.792 57.452 126.652 ;
    RECT 0.000 126.652 57.452 126.235 ;
    RECT 0.140 126.235 57.452 126.095 ;
    RECT 0.000 126.095 57.452 125.677 ;
    RECT 0.140 125.677 57.452 125.537 ;
    RECT 0.000 125.537 57.452 125.120 ;
    RECT 0.140 125.120 57.452 124.980 ;
    RECT 0.000 124.980 57.452 124.563 ;
    RECT 0.140 124.563 57.452 124.423 ;
    RECT 0.000 124.423 57.452 124.006 ;
    RECT 0.140 124.006 57.452 123.866 ;
    RECT 0.000 123.866 57.452 123.448 ;
    RECT 0.140 123.448 57.452 123.308 ;
    RECT 0.000 123.308 57.452 122.891 ;
    RECT 0.140 122.891 57.452 122.751 ;
    RECT 0.000 122.751 57.452 122.334 ;
    RECT 0.140 122.334 57.452 122.194 ;
    RECT 0.000 122.194 57.452 121.776 ;
    RECT 0.140 121.776 57.452 121.636 ;
    RECT 0.000 121.636 57.452 121.219 ;
    RECT 0.140 121.219 57.452 121.079 ;
    RECT 0.000 121.079 57.452 120.662 ;
    RECT 0.140 120.662 57.452 120.522 ;
    RECT 0.000 120.522 57.452 120.104 ;
    RECT 0.140 120.104 57.452 119.964 ;
    RECT 0.000 119.964 57.452 119.547 ;
    RECT 0.140 119.547 57.452 119.407 ;
    RECT 0.000 119.407 57.452 118.990 ;
    RECT 0.140 118.990 57.452 118.850 ;
    RECT 0.000 118.850 57.452 118.433 ;
    RECT 0.140 118.433 57.452 118.293 ;
    RECT 0.000 118.293 57.452 117.875 ;
    RECT 0.140 117.875 57.452 117.735 ;
    RECT 0.000 117.735 57.452 117.318 ;
    RECT 0.140 117.318 57.452 117.178 ;
    RECT 0.000 117.178 57.452 116.761 ;
    RECT 0.140 116.761 57.452 116.621 ;
    RECT 0.000 116.621 57.452 116.203 ;
    RECT 0.140 116.203 57.452 116.063 ;
    RECT 0.000 116.063 57.452 115.646 ;
    RECT 0.140 115.646 57.452 115.506 ;
    RECT 0.000 115.506 57.452 115.089 ;
    RECT 0.140 115.089 57.452 114.949 ;
    RECT 0.000 114.949 57.452 114.531 ;
    RECT 0.140 114.531 57.452 114.391 ;
    RECT 0.000 114.391 57.452 113.974 ;
    RECT 0.140 113.974 57.452 113.834 ;
    RECT 0.000 113.834 57.452 113.417 ;
    RECT 0.140 113.417 57.452 113.277 ;
    RECT 0.000 113.277 57.452 112.860 ;
    RECT 0.140 112.860 57.452 112.720 ;
    RECT 0.000 112.720 57.452 112.302 ;
    RECT 0.140 112.302 57.452 112.162 ;
    RECT 0.000 112.162 57.452 111.745 ;
    RECT 0.140 111.745 57.452 111.605 ;
    RECT 0.000 111.605 57.452 111.188 ;
    RECT 0.140 111.188 57.452 111.048 ;
    RECT 0.000 111.048 57.452 110.630 ;
    RECT 0.140 110.630 57.452 110.490 ;
    RECT 0.000 110.490 57.452 110.073 ;
    RECT 0.140 110.073 57.452 109.933 ;
    RECT 0.000 109.933 57.452 109.516 ;
    RECT 0.140 109.516 57.452 109.376 ;
    RECT 0.000 109.376 57.452 108.958 ;
    RECT 0.140 108.958 57.452 108.818 ;
    RECT 0.000 108.818 57.452 108.401 ;
    RECT 0.140 108.401 57.452 108.261 ;
    RECT 0.000 108.261 57.452 107.844 ;
    RECT 0.140 107.844 57.452 107.704 ;
    RECT 0.000 107.704 57.452 107.287 ;
    RECT 0.140 107.287 57.452 107.147 ;
    RECT 0.000 107.147 57.452 106.729 ;
    RECT 0.140 106.729 57.452 106.589 ;
    RECT 0.000 106.589 57.452 106.172 ;
    RECT 0.140 106.172 57.452 106.032 ;
    RECT 0.000 106.032 57.452 105.615 ;
    RECT 0.140 105.615 57.452 105.475 ;
    RECT 0.000 105.475 57.452 105.057 ;
    RECT 0.140 105.057 57.452 104.917 ;
    RECT 0.000 104.917 57.452 104.500 ;
    RECT 0.140 104.500 57.452 104.360 ;
    RECT 0.000 104.360 57.452 103.943 ;
    RECT 0.140 103.943 57.452 103.803 ;
    RECT 0.000 103.803 57.452 103.385 ;
    RECT 0.140 103.385 57.452 103.245 ;
    RECT 0.000 103.245 57.452 102.828 ;
    RECT 0.140 102.828 57.452 102.688 ;
    RECT 0.000 102.688 57.452 102.271 ;
    RECT 0.140 102.271 57.452 102.131 ;
    RECT 0.000 102.131 57.452 101.714 ;
    RECT 0.140 101.714 57.452 101.574 ;
    RECT 0.000 101.574 57.452 101.156 ;
    RECT 0.140 101.156 57.452 101.016 ;
    RECT 0.000 101.016 57.452 100.599 ;
    RECT 0.140 100.599 57.452 100.459 ;
    RECT 0.000 100.459 57.452 100.042 ;
    RECT 0.140 100.042 57.452 99.902 ;
    RECT 0.000 99.902 57.452 99.484 ;
    RECT 0.140 99.484 57.452 99.344 ;
    RECT 0.000 99.344 57.452 98.927 ;
    RECT 0.140 98.927 57.452 98.787 ;
    RECT 0.000 98.787 57.452 98.370 ;
    RECT 0.140 98.370 57.452 98.230 ;
    RECT 0.000 98.230 57.452 97.813 ;
    RECT 0.140 97.813 57.452 97.673 ;
    RECT 0.000 97.673 57.452 97.255 ;
    RECT 0.140 97.255 57.452 97.115 ;
    RECT 0.000 97.115 57.452 96.698 ;
    RECT 0.140 96.698 57.452 96.558 ;
    RECT 0.000 96.558 57.452 96.141 ;
    RECT 0.140 96.141 57.452 96.001 ;
    RECT 0.000 96.001 57.452 95.583 ;
    RECT 0.140 95.583 57.452 95.443 ;
    RECT 0.000 95.443 57.452 95.026 ;
    RECT 0.140 95.026 57.452 94.886 ;
    RECT 0.000 94.886 57.452 94.469 ;
    RECT 0.140 94.469 57.452 94.329 ;
    RECT 0.000 94.329 57.452 93.911 ;
    RECT 0.140 93.911 57.452 93.771 ;
    RECT 0.000 93.771 57.452 93.354 ;
    RECT 0.140 93.354 57.452 93.214 ;
    RECT 0.000 93.214 57.452 92.797 ;
    RECT 0.140 92.797 57.452 92.657 ;
    RECT 0.000 92.657 57.452 92.240 ;
    RECT 0.140 92.240 57.452 92.100 ;
    RECT 0.000 92.100 57.452 91.682 ;
    RECT 0.140 91.682 57.452 91.542 ;
    RECT 0.000 91.542 57.452 91.125 ;
    RECT 0.140 91.125 57.452 90.985 ;
    RECT 0.000 90.985 57.452 90.568 ;
    RECT 0.140 90.568 57.452 90.428 ;
    RECT 0.000 90.428 57.452 90.010 ;
    RECT 0.140 90.010 57.452 89.870 ;
    RECT 0.000 89.870 57.452 89.453 ;
    RECT 0.140 89.453 57.452 89.313 ;
    RECT 0.000 89.313 57.452 88.896 ;
    RECT 0.140 88.896 57.452 88.756 ;
    RECT 0.000 88.756 57.452 88.338 ;
    RECT 0.140 88.338 57.452 88.198 ;
    RECT 0.000 88.198 57.452 87.781 ;
    RECT 0.140 87.781 57.452 87.641 ;
    RECT 0.000 87.641 57.452 87.224 ;
    RECT 0.140 87.224 57.452 87.084 ;
    RECT 0.000 87.084 57.452 86.667 ;
    RECT 0.140 86.667 57.452 86.527 ;
    RECT 0.000 86.527 57.452 86.109 ;
    RECT 0.140 86.109 57.452 85.969 ;
    RECT 0.000 85.969 57.452 85.552 ;
    RECT 0.140 85.552 57.452 85.412 ;
    RECT 0.000 85.412 57.452 84.995 ;
    RECT 0.140 84.995 57.452 84.855 ;
    RECT 0.000 84.855 57.452 84.437 ;
    RECT 0.140 84.437 57.452 84.297 ;
    RECT 0.000 84.297 57.452 83.880 ;
    RECT 0.140 83.880 57.452 83.740 ;
    RECT 0.000 83.740 57.452 83.323 ;
    RECT 0.140 83.323 57.452 83.183 ;
    RECT 0.000 83.183 57.452 82.765 ;
    RECT 0.140 82.765 57.452 82.625 ;
    RECT 0.000 82.625 57.452 82.208 ;
    RECT 0.140 82.208 57.452 82.068 ;
    RECT 0.000 82.068 57.452 81.651 ;
    RECT 0.140 81.651 57.452 81.511 ;
    RECT 0.000 81.511 57.452 81.094 ;
    RECT 0.140 81.094 57.452 80.954 ;
    RECT 0.000 80.954 57.452 80.536 ;
    RECT 0.140 80.536 57.452 80.396 ;
    RECT 0.000 80.396 57.452 79.979 ;
    RECT 0.140 79.979 57.452 79.839 ;
    RECT 0.000 79.839 57.452 79.422 ;
    RECT 0.140 79.422 57.452 79.282 ;
    RECT 0.000 79.282 57.452 78.864 ;
    RECT 0.140 78.864 57.452 78.724 ;
    RECT 0.000 78.724 57.452 78.307 ;
    RECT 0.140 78.307 57.452 78.167 ;
    RECT 0.000 78.167 57.452 77.750 ;
    RECT 0.140 77.750 57.452 77.610 ;
    RECT 0.000 77.610 57.452 77.192 ;
    RECT 0.140 77.192 57.452 77.052 ;
    RECT 0.000 77.052 57.452 76.635 ;
    RECT 0.140 76.635 57.452 76.495 ;
    RECT 0.000 76.495 57.452 76.078 ;
    RECT 0.140 76.078 57.452 75.938 ;
    RECT 0.000 75.938 57.452 75.521 ;
    RECT 0.140 75.521 57.452 75.381 ;
    RECT 0.000 75.381 57.452 74.963 ;
    RECT 0.140 74.963 57.452 74.823 ;
    RECT 0.000 74.823 57.452 74.406 ;
    RECT 0.140 74.406 57.452 74.266 ;
    RECT 0.000 74.266 57.452 73.849 ;
    RECT 0.140 73.849 57.452 73.709 ;
    RECT 0.000 73.709 57.452 73.291 ;
    RECT 0.140 73.291 57.452 73.151 ;
    RECT 0.000 73.151 57.452 72.734 ;
    RECT 0.140 72.734 57.452 72.594 ;
    RECT 0.000 72.594 57.452 72.177 ;
    RECT 0.140 72.177 57.452 72.037 ;
    RECT 0.000 72.037 57.452 71.620 ;
    RECT 0.140 71.620 57.452 71.480 ;
    RECT 0.000 71.480 57.452 71.062 ;
    RECT 0.140 71.062 57.452 70.922 ;
    RECT 0.000 70.922 57.452 70.505 ;
    RECT 0.140 70.505 57.452 70.365 ;
    RECT 0.000 70.365 57.452 69.948 ;
    RECT 0.140 69.948 57.452 69.808 ;
    RECT 0.000 69.808 57.452 69.390 ;
    RECT 0.140 69.390 57.452 69.250 ;
    RECT 0.000 69.250 57.452 68.833 ;
    RECT 0.140 68.833 57.452 68.693 ;
    RECT 0.000 68.693 57.452 68.276 ;
    RECT 0.140 68.276 57.452 68.136 ;
    RECT 0.000 68.136 57.452 67.718 ;
    RECT 0.140 67.718 57.452 67.578 ;
    RECT 0.000 67.578 57.452 67.161 ;
    RECT 0.140 67.161 57.452 67.021 ;
    RECT 0.000 67.021 57.452 66.604 ;
    RECT 0.140 66.604 57.452 66.464 ;
    RECT 0.000 66.464 57.452 66.047 ;
    RECT 0.140 66.047 57.452 65.907 ;
    RECT 0.000 65.907 57.452 65.489 ;
    RECT 0.140 65.489 57.452 65.349 ;
    RECT 0.000 65.349 57.452 64.932 ;
    RECT 0.140 64.932 57.452 64.792 ;
    RECT 0.000 64.792 57.452 64.375 ;
    RECT 0.140 64.375 57.452 64.235 ;
    RECT 0.000 64.235 57.452 63.817 ;
    RECT 0.140 63.817 57.452 63.677 ;
    RECT 0.000 63.677 57.452 63.260 ;
    RECT 0.140 63.260 57.452 63.120 ;
    RECT 0.000 63.120 57.452 62.703 ;
    RECT 0.140 62.703 57.452 62.563 ;
    RECT 0.000 62.563 57.452 62.145 ;
    RECT 0.140 62.145 57.452 62.005 ;
    RECT 0.000 62.005 57.452 61.588 ;
    RECT 0.140 61.588 57.452 61.448 ;
    RECT 0.000 61.448 57.452 61.031 ;
    RECT 0.140 61.031 57.452 60.891 ;
    RECT 0.000 60.891 57.452 60.474 ;
    RECT 0.140 60.474 57.452 60.334 ;
    RECT 0.000 60.334 57.452 59.916 ;
    RECT 0.140 59.916 57.452 59.776 ;
    RECT 0.000 59.776 57.452 59.359 ;
    RECT 0.140 59.359 57.452 59.219 ;
    RECT 0.000 59.219 57.452 58.802 ;
    RECT 0.140 58.802 57.452 58.662 ;
    RECT 0.000 58.662 57.452 58.244 ;
    RECT 0.140 58.244 57.452 58.104 ;
    RECT 0.000 58.104 57.452 57.687 ;
    RECT 0.140 57.687 57.452 57.547 ;
    RECT 0.000 57.547 57.452 57.130 ;
    RECT 0.140 57.130 57.452 56.990 ;
    RECT 0.000 56.990 57.452 56.572 ;
    RECT 0.140 56.572 57.452 56.432 ;
    RECT 0.000 56.432 57.452 56.015 ;
    RECT 0.140 56.015 57.452 55.875 ;
    RECT 0.000 55.875 57.452 55.458 ;
    RECT 0.140 55.458 57.452 55.318 ;
    RECT 0.000 55.318 57.452 54.901 ;
    RECT 0.140 54.901 57.452 54.761 ;
    RECT 0.000 54.761 57.452 54.343 ;
    RECT 0.140 54.343 57.452 54.203 ;
    RECT 0.000 54.203 57.452 53.786 ;
    RECT 0.140 53.786 57.452 53.646 ;
    RECT 0.000 53.646 57.452 53.229 ;
    RECT 0.140 53.229 57.452 53.089 ;
    RECT 0.000 53.089 57.452 52.671 ;
    RECT 0.140 52.671 57.452 52.531 ;
    RECT 0.000 52.531 57.452 52.114 ;
    RECT 0.140 52.114 57.452 51.974 ;
    RECT 0.000 51.974 57.452 51.557 ;
    RECT 0.140 51.557 57.452 51.417 ;
    RECT 0.000 51.417 57.452 51.000 ;
    RECT 0.140 51.000 57.452 50.860 ;
    RECT 0.000 50.860 57.452 50.442 ;
    RECT 0.140 50.442 57.452 50.302 ;
    RECT 0.000 50.302 57.452 49.885 ;
    RECT 0.140 49.885 57.452 49.745 ;
    RECT 0.000 49.745 57.452 49.328 ;
    RECT 0.140 49.328 57.452 49.188 ;
    RECT 0.000 49.188 57.452 48.770 ;
    RECT 0.140 48.770 57.452 48.630 ;
    RECT 0.000 48.630 57.452 48.213 ;
    RECT 0.140 48.213 57.452 48.073 ;
    RECT 0.000 48.073 57.452 47.656 ;
    RECT 0.140 47.656 57.452 47.516 ;
    RECT 0.000 47.516 57.452 47.098 ;
    RECT 0.140 47.098 57.452 46.958 ;
    RECT 0.000 46.958 57.452 46.541 ;
    RECT 0.140 46.541 57.452 46.401 ;
    RECT 0.000 46.401 57.452 45.984 ;
    RECT 0.140 45.984 57.452 45.844 ;
    RECT 0.000 45.844 57.452 45.427 ;
    RECT 0.140 45.427 57.452 45.287 ;
    RECT 0.000 45.287 57.452 44.869 ;
    RECT 0.140 44.869 57.452 44.729 ;
    RECT 0.000 44.729 57.452 44.312 ;
    RECT 0.140 44.312 57.452 44.172 ;
    RECT 0.000 44.172 57.452 43.755 ;
    RECT 0.140 43.755 57.452 43.615 ;
    RECT 0.000 43.615 57.452 43.197 ;
    RECT 0.140 43.197 57.452 43.057 ;
    RECT 0.000 43.057 57.452 42.640 ;
    RECT 0.140 42.640 57.452 42.500 ;
    RECT 0.000 42.500 57.452 42.083 ;
    RECT 0.140 42.083 57.452 41.943 ;
    RECT 0.000 41.943 57.452 41.525 ;
    RECT 0.140 41.525 57.452 41.385 ;
    RECT 0.000 41.385 57.452 40.968 ;
    RECT 0.140 40.968 57.452 40.828 ;
    RECT 0.000 40.828 57.452 40.411 ;
    RECT 0.140 40.411 57.452 40.271 ;
    RECT 0.000 40.271 57.452 39.854 ;
    RECT 0.140 39.854 57.452 39.714 ;
    RECT 0.000 39.714 57.452 39.296 ;
    RECT 0.140 39.296 57.452 39.156 ;
    RECT 0.000 39.156 57.452 38.739 ;
    RECT 0.140 38.739 57.452 38.599 ;
    RECT 0.000 38.599 57.452 38.182 ;
    RECT 0.140 38.182 57.452 38.042 ;
    RECT 0.000 38.042 57.452 37.624 ;
    RECT 0.140 37.624 57.452 37.484 ;
    RECT 0.000 37.484 57.452 37.067 ;
    RECT 0.140 37.067 57.452 36.927 ;
    RECT 0.000 36.927 57.452 36.510 ;
    RECT 0.140 36.510 57.452 36.370 ;
    RECT 0.000 36.370 57.452 35.952 ;
    RECT 0.140 35.952 57.452 35.812 ;
    RECT 0.000 35.812 57.452 35.395 ;
    RECT 0.140 35.395 57.452 35.255 ;
    RECT 0.000 35.255 57.452 34.838 ;
    RECT 0.140 34.838 57.452 34.698 ;
    RECT 0.000 34.698 57.452 34.281 ;
    RECT 0.140 34.281 57.452 34.141 ;
    RECT 0.000 34.141 57.452 33.723 ;
    RECT 0.140 33.723 57.452 33.583 ;
    RECT 0.000 33.583 57.452 33.166 ;
    RECT 0.140 33.166 57.452 33.026 ;
    RECT 0.000 33.026 57.452 32.609 ;
    RECT 0.140 32.609 57.452 32.469 ;
    RECT 0.000 32.469 57.452 32.051 ;
    RECT 0.140 32.051 57.452 31.911 ;
    RECT 0.000 31.911 57.452 31.494 ;
    RECT 0.140 31.494 57.452 31.354 ;
    RECT 0.000 31.354 57.452 30.937 ;
    RECT 0.140 30.937 57.452 30.797 ;
    RECT 0.000 30.797 57.452 30.379 ;
    RECT 0.140 30.379 57.452 30.239 ;
    RECT 0.000 30.239 57.452 29.822 ;
    RECT 0.140 29.822 57.452 29.682 ;
    RECT 0.000 29.682 57.452 29.265 ;
    RECT 0.140 29.265 57.452 29.125 ;
    RECT 0.000 29.125 57.452 28.708 ;
    RECT 0.140 28.708 57.452 28.568 ;
    RECT 0.000 28.568 57.452 28.150 ;
    RECT 0.140 28.150 57.452 28.010 ;
    RECT 0.000 28.010 57.452 27.593 ;
    RECT 0.140 27.593 57.452 27.453 ;
    RECT 0.000 27.453 57.452 27.036 ;
    RECT 0.140 27.036 57.452 26.896 ;
    RECT 0.000 26.896 57.452 26.478 ;
    RECT 0.140 26.478 57.452 26.338 ;
    RECT 0.000 26.338 57.452 25.921 ;
    RECT 0.140 25.921 57.452 25.781 ;
    RECT 0.000 25.781 57.452 25.364 ;
    RECT 0.140 25.364 57.452 25.224 ;
    RECT 0.000 25.224 57.452 24.807 ;
    RECT 0.140 24.807 57.452 24.667 ;
    RECT 0.000 24.667 57.452 24.249 ;
    RECT 0.140 24.249 57.452 24.109 ;
    RECT 0.000 24.109 57.452 23.692 ;
    RECT 0.140 23.692 57.452 23.552 ;
    RECT 0.000 23.552 57.452 23.135 ;
    RECT 0.140 23.135 57.452 22.995 ;
    RECT 0.000 22.995 57.452 22.577 ;
    RECT 0.140 22.577 57.452 22.437 ;
    RECT 0.000 22.437 57.452 22.020 ;
    RECT 0.140 22.020 57.452 21.880 ;
    RECT 0.000 21.880 57.452 21.463 ;
    RECT 0.140 21.463 57.452 21.323 ;
    RECT 0.000 21.323 57.452 20.905 ;
    RECT 0.140 20.905 57.452 20.765 ;
    RECT 0.000 20.765 57.452 20.348 ;
    RECT 0.140 20.348 57.452 20.208 ;
    RECT 0.000 20.208 57.452 19.791 ;
    RECT 0.140 19.791 57.452 19.651 ;
    RECT 0.000 19.651 57.452 19.234 ;
    RECT 0.140 19.234 57.452 19.094 ;
    RECT 0.000 19.094 57.452 18.676 ;
    RECT 0.140 18.676 57.452 18.536 ;
    RECT 0.000 18.536 57.452 18.119 ;
    RECT 0.140 18.119 57.452 17.979 ;
    RECT 0.000 17.979 57.452 17.562 ;
    RECT 0.140 17.562 57.452 17.422 ;
    RECT 0.000 17.422 57.452 17.004 ;
    RECT 0.140 17.004 57.452 16.864 ;
    RECT 0.000 16.864 57.452 16.447 ;
    RECT 0.140 16.447 57.452 16.307 ;
    RECT 0.000 16.307 57.452 15.890 ;
    RECT 0.140 15.890 57.452 15.750 ;
    RECT 0.000 15.750 57.452 15.332 ;
    RECT 0.140 15.332 57.452 15.192 ;
    RECT 0.000 15.192 57.452 14.775 ;
    RECT 0.140 14.775 57.452 14.635 ;
    RECT 0.000 14.635 57.452 14.218 ;
    RECT 0.140 14.218 57.452 14.078 ;
    RECT 0.000 14.078 57.452 13.661 ;
    RECT 0.140 13.661 57.452 13.521 ;
    RECT 0.000 13.521 57.452 13.103 ;
    RECT 0.140 13.103 57.452 12.963 ;
    RECT 0.000 12.963 57.452 12.546 ;
    RECT 0.140 12.546 57.452 12.406 ;
    RECT 0.000 12.406 57.452 11.989 ;
    RECT 0.140 11.989 57.452 11.849 ;
    RECT 0.000 11.849 57.452 11.431 ;
    RECT 0.140 11.431 57.452 11.291 ;
    RECT 0.000 11.291 57.452 10.874 ;
    RECT 0.140 10.874 57.452 10.734 ;
    RECT 0.000 10.734 57.452 10.317 ;
    RECT 0.140 10.317 57.452 10.177 ;
    RECT 0.000 10.177 57.452 9.759 ;
    RECT 0.140 9.759 57.452 9.619 ;
    RECT 0.000 9.619 57.452 9.202 ;
    RECT 0.140 9.202 57.452 9.062 ;
    RECT 0.000 9.062 57.452 8.645 ;
    RECT 0.140 8.645 57.452 8.505 ;
    RECT 0.000 8.505 57.452 8.088 ;
    RECT 0.140 8.088 57.452 7.948 ;
    RECT 0.000 7.948 57.452 7.530 ;
    RECT 0.140 7.530 57.452 7.390 ;
    RECT 0.000 7.390 57.452 6.973 ;
    RECT 0.140 6.973 57.452 6.833 ;
    RECT 0.000 6.833 57.452 6.416 ;
    RECT 0.140 6.416 57.452 6.276 ;
    RECT 0.000 6.276 57.452 5.858 ;
    RECT 0.140 5.858 57.452 5.718 ;
    RECT 0.000 5.718 57.452 5.301 ;
    RECT 0.140 5.301 57.452 5.161 ;
    RECT 0.000 5.161 57.452 4.744 ;
    RECT 0.140 4.744 57.452 4.604 ;
    RECT 0.000 4.604 57.452 4.186 ;
    RECT 0.140 4.186 57.452 4.046 ;
    RECT 0.000 4.046 57.452 3.629 ;
    RECT 0.140 3.629 57.452 3.489 ;
    RECT 0.000 3.489 57.452 3.072 ;
    RECT 0.140 3.072 57.452 2.932 ;
    RECT 0.000 2.932 57.452 2.515 ;
    RECT 0.140 2.515 57.452 2.375 ;
    RECT 0.000 2.375 57.452 1.957 ;
    RECT 0.140 1.957 57.452 1.817 ;
    RECT 0.000 1.817 57.452 1.400 ;
    RECT 0.000 1.400 57.452 0.000 ;
    LAYER metal3 ;
    RECT 0.000 167.760 57.452 166.360 ;
    RECT 0.140 166.360 57.452 166.220 ;
    RECT 0.000 166.220 57.452 165.803 ;
    RECT 0.140 165.803 57.452 165.663 ;
    RECT 0.000 165.663 57.452 165.246 ;
    RECT 0.140 165.246 57.452 165.106 ;
    RECT 0.000 165.106 57.452 164.688 ;
    RECT 0.140 164.688 57.452 164.548 ;
    RECT 0.000 164.548 57.452 164.131 ;
    RECT 0.140 164.131 57.452 163.991 ;
    RECT 0.000 163.991 57.452 163.574 ;
    RECT 0.140 163.574 57.452 163.434 ;
    RECT 0.000 163.434 57.452 163.016 ;
    RECT 0.140 163.016 57.452 162.876 ;
    RECT 0.000 162.876 57.452 162.459 ;
    RECT 0.140 162.459 57.452 162.319 ;
    RECT 0.000 162.319 57.452 161.902 ;
    RECT 0.140 161.902 57.452 161.762 ;
    RECT 0.000 161.762 57.452 161.344 ;
    RECT 0.140 161.344 57.452 161.204 ;
    RECT 0.000 161.204 57.452 160.787 ;
    RECT 0.140 160.787 57.452 160.647 ;
    RECT 0.000 160.647 57.452 160.230 ;
    RECT 0.140 160.230 57.452 160.090 ;
    RECT 0.000 160.090 57.452 159.673 ;
    RECT 0.140 159.673 57.452 159.533 ;
    RECT 0.000 159.533 57.452 159.115 ;
    RECT 0.140 159.115 57.452 158.975 ;
    RECT 0.000 158.975 57.452 158.558 ;
    RECT 0.140 158.558 57.452 158.418 ;
    RECT 0.000 158.418 57.452 158.001 ;
    RECT 0.140 158.001 57.452 157.861 ;
    RECT 0.000 157.861 57.452 157.443 ;
    RECT 0.140 157.443 57.452 157.303 ;
    RECT 0.000 157.303 57.452 156.886 ;
    RECT 0.140 156.886 57.452 156.746 ;
    RECT 0.000 156.746 57.452 156.329 ;
    RECT 0.140 156.329 57.452 156.189 ;
    RECT 0.000 156.189 57.452 155.771 ;
    RECT 0.140 155.771 57.452 155.631 ;
    RECT 0.000 155.631 57.452 155.214 ;
    RECT 0.140 155.214 57.452 155.074 ;
    RECT 0.000 155.074 57.452 154.657 ;
    RECT 0.140 154.657 57.452 154.517 ;
    RECT 0.000 154.517 57.452 154.100 ;
    RECT 0.140 154.100 57.452 153.960 ;
    RECT 0.000 153.960 57.452 153.542 ;
    RECT 0.140 153.542 57.452 153.402 ;
    RECT 0.000 153.402 57.452 152.985 ;
    RECT 0.140 152.985 57.452 152.845 ;
    RECT 0.000 152.845 57.452 152.428 ;
    RECT 0.140 152.428 57.452 152.288 ;
    RECT 0.000 152.288 57.452 151.870 ;
    RECT 0.140 151.870 57.452 151.730 ;
    RECT 0.000 151.730 57.452 151.313 ;
    RECT 0.140 151.313 57.452 151.173 ;
    RECT 0.000 151.173 57.452 150.756 ;
    RECT 0.140 150.756 57.452 150.616 ;
    RECT 0.000 150.616 57.452 150.199 ;
    RECT 0.140 150.199 57.452 150.059 ;
    RECT 0.000 150.059 57.452 149.641 ;
    RECT 0.140 149.641 57.452 149.501 ;
    RECT 0.000 149.501 57.452 149.084 ;
    RECT 0.140 149.084 57.452 148.944 ;
    RECT 0.000 148.944 57.452 148.527 ;
    RECT 0.140 148.527 57.452 148.387 ;
    RECT 0.000 148.387 57.452 147.969 ;
    RECT 0.140 147.969 57.452 147.829 ;
    RECT 0.000 147.829 57.452 147.412 ;
    RECT 0.140 147.412 57.452 147.272 ;
    RECT 0.000 147.272 57.452 146.855 ;
    RECT 0.140 146.855 57.452 146.715 ;
    RECT 0.000 146.715 57.452 146.297 ;
    RECT 0.140 146.297 57.452 146.157 ;
    RECT 0.000 146.157 57.452 145.740 ;
    RECT 0.140 145.740 57.452 145.600 ;
    RECT 0.000 145.600 57.452 145.183 ;
    RECT 0.140 145.183 57.452 145.043 ;
    RECT 0.000 145.043 57.452 144.626 ;
    RECT 0.140 144.626 57.452 144.486 ;
    RECT 0.000 144.486 57.452 144.068 ;
    RECT 0.140 144.068 57.452 143.928 ;
    RECT 0.000 143.928 57.452 143.511 ;
    RECT 0.140 143.511 57.452 143.371 ;
    RECT 0.000 143.371 57.452 142.954 ;
    RECT 0.140 142.954 57.452 142.814 ;
    RECT 0.000 142.814 57.452 142.396 ;
    RECT 0.140 142.396 57.452 142.256 ;
    RECT 0.000 142.256 57.452 141.839 ;
    RECT 0.140 141.839 57.452 141.699 ;
    RECT 0.000 141.699 57.452 141.282 ;
    RECT 0.140 141.282 57.452 141.142 ;
    RECT 0.000 141.142 57.452 140.724 ;
    RECT 0.140 140.724 57.452 140.584 ;
    RECT 0.000 140.584 57.452 140.167 ;
    RECT 0.140 140.167 57.452 140.027 ;
    RECT 0.000 140.027 57.452 139.610 ;
    RECT 0.140 139.610 57.452 139.470 ;
    RECT 0.000 139.470 57.452 139.053 ;
    RECT 0.140 139.053 57.452 138.913 ;
    RECT 0.000 138.913 57.452 138.495 ;
    RECT 0.140 138.495 57.452 138.355 ;
    RECT 0.000 138.355 57.452 137.938 ;
    RECT 0.140 137.938 57.452 137.798 ;
    RECT 0.000 137.798 57.452 137.381 ;
    RECT 0.140 137.381 57.452 137.241 ;
    RECT 0.000 137.241 57.452 136.823 ;
    RECT 0.140 136.823 57.452 136.683 ;
    RECT 0.000 136.683 57.452 136.266 ;
    RECT 0.140 136.266 57.452 136.126 ;
    RECT 0.000 136.126 57.452 135.709 ;
    RECT 0.140 135.709 57.452 135.569 ;
    RECT 0.000 135.569 57.452 135.151 ;
    RECT 0.140 135.151 57.452 135.011 ;
    RECT 0.000 135.011 57.452 134.594 ;
    RECT 0.140 134.594 57.452 134.454 ;
    RECT 0.000 134.454 57.452 134.037 ;
    RECT 0.140 134.037 57.452 133.897 ;
    RECT 0.000 133.897 57.452 133.480 ;
    RECT 0.140 133.480 57.452 133.340 ;
    RECT 0.000 133.340 57.452 132.922 ;
    RECT 0.140 132.922 57.452 132.782 ;
    RECT 0.000 132.782 57.452 132.365 ;
    RECT 0.140 132.365 57.452 132.225 ;
    RECT 0.000 132.225 57.452 131.808 ;
    RECT 0.140 131.808 57.452 131.668 ;
    RECT 0.000 131.668 57.452 131.250 ;
    RECT 0.140 131.250 57.452 131.110 ;
    RECT 0.000 131.110 57.452 130.693 ;
    RECT 0.140 130.693 57.452 130.553 ;
    RECT 0.000 130.553 57.452 130.136 ;
    RECT 0.140 130.136 57.452 129.996 ;
    RECT 0.000 129.996 57.452 129.578 ;
    RECT 0.140 129.578 57.452 129.438 ;
    RECT 0.000 129.438 57.452 129.021 ;
    RECT 0.140 129.021 57.452 128.881 ;
    RECT 0.000 128.881 57.452 128.464 ;
    RECT 0.140 128.464 57.452 128.324 ;
    RECT 0.000 128.324 57.452 127.907 ;
    RECT 0.140 127.907 57.452 127.767 ;
    RECT 0.000 127.767 57.452 127.349 ;
    RECT 0.140 127.349 57.452 127.209 ;
    RECT 0.000 127.209 57.452 126.792 ;
    RECT 0.140 126.792 57.452 126.652 ;
    RECT 0.000 126.652 57.452 126.235 ;
    RECT 0.140 126.235 57.452 126.095 ;
    RECT 0.000 126.095 57.452 125.677 ;
    RECT 0.140 125.677 57.452 125.537 ;
    RECT 0.000 125.537 57.452 125.120 ;
    RECT 0.140 125.120 57.452 124.980 ;
    RECT 0.000 124.980 57.452 124.563 ;
    RECT 0.140 124.563 57.452 124.423 ;
    RECT 0.000 124.423 57.452 124.006 ;
    RECT 0.140 124.006 57.452 123.866 ;
    RECT 0.000 123.866 57.452 123.448 ;
    RECT 0.140 123.448 57.452 123.308 ;
    RECT 0.000 123.308 57.452 122.891 ;
    RECT 0.140 122.891 57.452 122.751 ;
    RECT 0.000 122.751 57.452 122.334 ;
    RECT 0.140 122.334 57.452 122.194 ;
    RECT 0.000 122.194 57.452 121.776 ;
    RECT 0.140 121.776 57.452 121.636 ;
    RECT 0.000 121.636 57.452 121.219 ;
    RECT 0.140 121.219 57.452 121.079 ;
    RECT 0.000 121.079 57.452 120.662 ;
    RECT 0.140 120.662 57.452 120.522 ;
    RECT 0.000 120.522 57.452 120.104 ;
    RECT 0.140 120.104 57.452 119.964 ;
    RECT 0.000 119.964 57.452 119.547 ;
    RECT 0.140 119.547 57.452 119.407 ;
    RECT 0.000 119.407 57.452 118.990 ;
    RECT 0.140 118.990 57.452 118.850 ;
    RECT 0.000 118.850 57.452 118.433 ;
    RECT 0.140 118.433 57.452 118.293 ;
    RECT 0.000 118.293 57.452 117.875 ;
    RECT 0.140 117.875 57.452 117.735 ;
    RECT 0.000 117.735 57.452 117.318 ;
    RECT 0.140 117.318 57.452 117.178 ;
    RECT 0.000 117.178 57.452 116.761 ;
    RECT 0.140 116.761 57.452 116.621 ;
    RECT 0.000 116.621 57.452 116.203 ;
    RECT 0.140 116.203 57.452 116.063 ;
    RECT 0.000 116.063 57.452 115.646 ;
    RECT 0.140 115.646 57.452 115.506 ;
    RECT 0.000 115.506 57.452 115.089 ;
    RECT 0.140 115.089 57.452 114.949 ;
    RECT 0.000 114.949 57.452 114.531 ;
    RECT 0.140 114.531 57.452 114.391 ;
    RECT 0.000 114.391 57.452 113.974 ;
    RECT 0.140 113.974 57.452 113.834 ;
    RECT 0.000 113.834 57.452 113.417 ;
    RECT 0.140 113.417 57.452 113.277 ;
    RECT 0.000 113.277 57.452 112.860 ;
    RECT 0.140 112.860 57.452 112.720 ;
    RECT 0.000 112.720 57.452 112.302 ;
    RECT 0.140 112.302 57.452 112.162 ;
    RECT 0.000 112.162 57.452 111.745 ;
    RECT 0.140 111.745 57.452 111.605 ;
    RECT 0.000 111.605 57.452 111.188 ;
    RECT 0.140 111.188 57.452 111.048 ;
    RECT 0.000 111.048 57.452 110.630 ;
    RECT 0.140 110.630 57.452 110.490 ;
    RECT 0.000 110.490 57.452 110.073 ;
    RECT 0.140 110.073 57.452 109.933 ;
    RECT 0.000 109.933 57.452 109.516 ;
    RECT 0.140 109.516 57.452 109.376 ;
    RECT 0.000 109.376 57.452 108.958 ;
    RECT 0.140 108.958 57.452 108.818 ;
    RECT 0.000 108.818 57.452 108.401 ;
    RECT 0.140 108.401 57.452 108.261 ;
    RECT 0.000 108.261 57.452 107.844 ;
    RECT 0.140 107.844 57.452 107.704 ;
    RECT 0.000 107.704 57.452 107.287 ;
    RECT 0.140 107.287 57.452 107.147 ;
    RECT 0.000 107.147 57.452 106.729 ;
    RECT 0.140 106.729 57.452 106.589 ;
    RECT 0.000 106.589 57.452 106.172 ;
    RECT 0.140 106.172 57.452 106.032 ;
    RECT 0.000 106.032 57.452 105.615 ;
    RECT 0.140 105.615 57.452 105.475 ;
    RECT 0.000 105.475 57.452 105.057 ;
    RECT 0.140 105.057 57.452 104.917 ;
    RECT 0.000 104.917 57.452 104.500 ;
    RECT 0.140 104.500 57.452 104.360 ;
    RECT 0.000 104.360 57.452 103.943 ;
    RECT 0.140 103.943 57.452 103.803 ;
    RECT 0.000 103.803 57.452 103.385 ;
    RECT 0.140 103.385 57.452 103.245 ;
    RECT 0.000 103.245 57.452 102.828 ;
    RECT 0.140 102.828 57.452 102.688 ;
    RECT 0.000 102.688 57.452 102.271 ;
    RECT 0.140 102.271 57.452 102.131 ;
    RECT 0.000 102.131 57.452 101.714 ;
    RECT 0.140 101.714 57.452 101.574 ;
    RECT 0.000 101.574 57.452 101.156 ;
    RECT 0.140 101.156 57.452 101.016 ;
    RECT 0.000 101.016 57.452 100.599 ;
    RECT 0.140 100.599 57.452 100.459 ;
    RECT 0.000 100.459 57.452 100.042 ;
    RECT 0.140 100.042 57.452 99.902 ;
    RECT 0.000 99.902 57.452 99.484 ;
    RECT 0.140 99.484 57.452 99.344 ;
    RECT 0.000 99.344 57.452 98.927 ;
    RECT 0.140 98.927 57.452 98.787 ;
    RECT 0.000 98.787 57.452 98.370 ;
    RECT 0.140 98.370 57.452 98.230 ;
    RECT 0.000 98.230 57.452 97.813 ;
    RECT 0.140 97.813 57.452 97.673 ;
    RECT 0.000 97.673 57.452 97.255 ;
    RECT 0.140 97.255 57.452 97.115 ;
    RECT 0.000 97.115 57.452 96.698 ;
    RECT 0.140 96.698 57.452 96.558 ;
    RECT 0.000 96.558 57.452 96.141 ;
    RECT 0.140 96.141 57.452 96.001 ;
    RECT 0.000 96.001 57.452 95.583 ;
    RECT 0.140 95.583 57.452 95.443 ;
    RECT 0.000 95.443 57.452 95.026 ;
    RECT 0.140 95.026 57.452 94.886 ;
    RECT 0.000 94.886 57.452 94.469 ;
    RECT 0.140 94.469 57.452 94.329 ;
    RECT 0.000 94.329 57.452 93.911 ;
    RECT 0.140 93.911 57.452 93.771 ;
    RECT 0.000 93.771 57.452 93.354 ;
    RECT 0.140 93.354 57.452 93.214 ;
    RECT 0.000 93.214 57.452 92.797 ;
    RECT 0.140 92.797 57.452 92.657 ;
    RECT 0.000 92.657 57.452 92.240 ;
    RECT 0.140 92.240 57.452 92.100 ;
    RECT 0.000 92.100 57.452 91.682 ;
    RECT 0.140 91.682 57.452 91.542 ;
    RECT 0.000 91.542 57.452 91.125 ;
    RECT 0.140 91.125 57.452 90.985 ;
    RECT 0.000 90.985 57.452 90.568 ;
    RECT 0.140 90.568 57.452 90.428 ;
    RECT 0.000 90.428 57.452 90.010 ;
    RECT 0.140 90.010 57.452 89.870 ;
    RECT 0.000 89.870 57.452 89.453 ;
    RECT 0.140 89.453 57.452 89.313 ;
    RECT 0.000 89.313 57.452 88.896 ;
    RECT 0.140 88.896 57.452 88.756 ;
    RECT 0.000 88.756 57.452 88.338 ;
    RECT 0.140 88.338 57.452 88.198 ;
    RECT 0.000 88.198 57.452 87.781 ;
    RECT 0.140 87.781 57.452 87.641 ;
    RECT 0.000 87.641 57.452 87.224 ;
    RECT 0.140 87.224 57.452 87.084 ;
    RECT 0.000 87.084 57.452 86.667 ;
    RECT 0.140 86.667 57.452 86.527 ;
    RECT 0.000 86.527 57.452 86.109 ;
    RECT 0.140 86.109 57.452 85.969 ;
    RECT 0.000 85.969 57.452 85.552 ;
    RECT 0.140 85.552 57.452 85.412 ;
    RECT 0.000 85.412 57.452 84.995 ;
    RECT 0.140 84.995 57.452 84.855 ;
    RECT 0.000 84.855 57.452 84.437 ;
    RECT 0.140 84.437 57.452 84.297 ;
    RECT 0.000 84.297 57.452 83.880 ;
    RECT 0.140 83.880 57.452 83.740 ;
    RECT 0.000 83.740 57.452 83.323 ;
    RECT 0.140 83.323 57.452 83.183 ;
    RECT 0.000 83.183 57.452 82.765 ;
    RECT 0.140 82.765 57.452 82.625 ;
    RECT 0.000 82.625 57.452 82.208 ;
    RECT 0.140 82.208 57.452 82.068 ;
    RECT 0.000 82.068 57.452 81.651 ;
    RECT 0.140 81.651 57.452 81.511 ;
    RECT 0.000 81.511 57.452 81.094 ;
    RECT 0.140 81.094 57.452 80.954 ;
    RECT 0.000 80.954 57.452 80.536 ;
    RECT 0.140 80.536 57.452 80.396 ;
    RECT 0.000 80.396 57.452 79.979 ;
    RECT 0.140 79.979 57.452 79.839 ;
    RECT 0.000 79.839 57.452 79.422 ;
    RECT 0.140 79.422 57.452 79.282 ;
    RECT 0.000 79.282 57.452 78.864 ;
    RECT 0.140 78.864 57.452 78.724 ;
    RECT 0.000 78.724 57.452 78.307 ;
    RECT 0.140 78.307 57.452 78.167 ;
    RECT 0.000 78.167 57.452 77.750 ;
    RECT 0.140 77.750 57.452 77.610 ;
    RECT 0.000 77.610 57.452 77.192 ;
    RECT 0.140 77.192 57.452 77.052 ;
    RECT 0.000 77.052 57.452 76.635 ;
    RECT 0.140 76.635 57.452 76.495 ;
    RECT 0.000 76.495 57.452 76.078 ;
    RECT 0.140 76.078 57.452 75.938 ;
    RECT 0.000 75.938 57.452 75.521 ;
    RECT 0.140 75.521 57.452 75.381 ;
    RECT 0.000 75.381 57.452 74.963 ;
    RECT 0.140 74.963 57.452 74.823 ;
    RECT 0.000 74.823 57.452 74.406 ;
    RECT 0.140 74.406 57.452 74.266 ;
    RECT 0.000 74.266 57.452 73.849 ;
    RECT 0.140 73.849 57.452 73.709 ;
    RECT 0.000 73.709 57.452 73.291 ;
    RECT 0.140 73.291 57.452 73.151 ;
    RECT 0.000 73.151 57.452 72.734 ;
    RECT 0.140 72.734 57.452 72.594 ;
    RECT 0.000 72.594 57.452 72.177 ;
    RECT 0.140 72.177 57.452 72.037 ;
    RECT 0.000 72.037 57.452 71.620 ;
    RECT 0.140 71.620 57.452 71.480 ;
    RECT 0.000 71.480 57.452 71.062 ;
    RECT 0.140 71.062 57.452 70.922 ;
    RECT 0.000 70.922 57.452 70.505 ;
    RECT 0.140 70.505 57.452 70.365 ;
    RECT 0.000 70.365 57.452 69.948 ;
    RECT 0.140 69.948 57.452 69.808 ;
    RECT 0.000 69.808 57.452 69.390 ;
    RECT 0.140 69.390 57.452 69.250 ;
    RECT 0.000 69.250 57.452 68.833 ;
    RECT 0.140 68.833 57.452 68.693 ;
    RECT 0.000 68.693 57.452 68.276 ;
    RECT 0.140 68.276 57.452 68.136 ;
    RECT 0.000 68.136 57.452 67.718 ;
    RECT 0.140 67.718 57.452 67.578 ;
    RECT 0.000 67.578 57.452 67.161 ;
    RECT 0.140 67.161 57.452 67.021 ;
    RECT 0.000 67.021 57.452 66.604 ;
    RECT 0.140 66.604 57.452 66.464 ;
    RECT 0.000 66.464 57.452 66.047 ;
    RECT 0.140 66.047 57.452 65.907 ;
    RECT 0.000 65.907 57.452 65.489 ;
    RECT 0.140 65.489 57.452 65.349 ;
    RECT 0.000 65.349 57.452 64.932 ;
    RECT 0.140 64.932 57.452 64.792 ;
    RECT 0.000 64.792 57.452 64.375 ;
    RECT 0.140 64.375 57.452 64.235 ;
    RECT 0.000 64.235 57.452 63.817 ;
    RECT 0.140 63.817 57.452 63.677 ;
    RECT 0.000 63.677 57.452 63.260 ;
    RECT 0.140 63.260 57.452 63.120 ;
    RECT 0.000 63.120 57.452 62.703 ;
    RECT 0.140 62.703 57.452 62.563 ;
    RECT 0.000 62.563 57.452 62.145 ;
    RECT 0.140 62.145 57.452 62.005 ;
    RECT 0.000 62.005 57.452 61.588 ;
    RECT 0.140 61.588 57.452 61.448 ;
    RECT 0.000 61.448 57.452 61.031 ;
    RECT 0.140 61.031 57.452 60.891 ;
    RECT 0.000 60.891 57.452 60.474 ;
    RECT 0.140 60.474 57.452 60.334 ;
    RECT 0.000 60.334 57.452 59.916 ;
    RECT 0.140 59.916 57.452 59.776 ;
    RECT 0.000 59.776 57.452 59.359 ;
    RECT 0.140 59.359 57.452 59.219 ;
    RECT 0.000 59.219 57.452 58.802 ;
    RECT 0.140 58.802 57.452 58.662 ;
    RECT 0.000 58.662 57.452 58.244 ;
    RECT 0.140 58.244 57.452 58.104 ;
    RECT 0.000 58.104 57.452 57.687 ;
    RECT 0.140 57.687 57.452 57.547 ;
    RECT 0.000 57.547 57.452 57.130 ;
    RECT 0.140 57.130 57.452 56.990 ;
    RECT 0.000 56.990 57.452 56.572 ;
    RECT 0.140 56.572 57.452 56.432 ;
    RECT 0.000 56.432 57.452 56.015 ;
    RECT 0.140 56.015 57.452 55.875 ;
    RECT 0.000 55.875 57.452 55.458 ;
    RECT 0.140 55.458 57.452 55.318 ;
    RECT 0.000 55.318 57.452 54.901 ;
    RECT 0.140 54.901 57.452 54.761 ;
    RECT 0.000 54.761 57.452 54.343 ;
    RECT 0.140 54.343 57.452 54.203 ;
    RECT 0.000 54.203 57.452 53.786 ;
    RECT 0.140 53.786 57.452 53.646 ;
    RECT 0.000 53.646 57.452 53.229 ;
    RECT 0.140 53.229 57.452 53.089 ;
    RECT 0.000 53.089 57.452 52.671 ;
    RECT 0.140 52.671 57.452 52.531 ;
    RECT 0.000 52.531 57.452 52.114 ;
    RECT 0.140 52.114 57.452 51.974 ;
    RECT 0.000 51.974 57.452 51.557 ;
    RECT 0.140 51.557 57.452 51.417 ;
    RECT 0.000 51.417 57.452 51.000 ;
    RECT 0.140 51.000 57.452 50.860 ;
    RECT 0.000 50.860 57.452 50.442 ;
    RECT 0.140 50.442 57.452 50.302 ;
    RECT 0.000 50.302 57.452 49.885 ;
    RECT 0.140 49.885 57.452 49.745 ;
    RECT 0.000 49.745 57.452 49.328 ;
    RECT 0.140 49.328 57.452 49.188 ;
    RECT 0.000 49.188 57.452 48.770 ;
    RECT 0.140 48.770 57.452 48.630 ;
    RECT 0.000 48.630 57.452 48.213 ;
    RECT 0.140 48.213 57.452 48.073 ;
    RECT 0.000 48.073 57.452 47.656 ;
    RECT 0.140 47.656 57.452 47.516 ;
    RECT 0.000 47.516 57.452 47.098 ;
    RECT 0.140 47.098 57.452 46.958 ;
    RECT 0.000 46.958 57.452 46.541 ;
    RECT 0.140 46.541 57.452 46.401 ;
    RECT 0.000 46.401 57.452 45.984 ;
    RECT 0.140 45.984 57.452 45.844 ;
    RECT 0.000 45.844 57.452 45.427 ;
    RECT 0.140 45.427 57.452 45.287 ;
    RECT 0.000 45.287 57.452 44.869 ;
    RECT 0.140 44.869 57.452 44.729 ;
    RECT 0.000 44.729 57.452 44.312 ;
    RECT 0.140 44.312 57.452 44.172 ;
    RECT 0.000 44.172 57.452 43.755 ;
    RECT 0.140 43.755 57.452 43.615 ;
    RECT 0.000 43.615 57.452 43.197 ;
    RECT 0.140 43.197 57.452 43.057 ;
    RECT 0.000 43.057 57.452 42.640 ;
    RECT 0.140 42.640 57.452 42.500 ;
    RECT 0.000 42.500 57.452 42.083 ;
    RECT 0.140 42.083 57.452 41.943 ;
    RECT 0.000 41.943 57.452 41.525 ;
    RECT 0.140 41.525 57.452 41.385 ;
    RECT 0.000 41.385 57.452 40.968 ;
    RECT 0.140 40.968 57.452 40.828 ;
    RECT 0.000 40.828 57.452 40.411 ;
    RECT 0.140 40.411 57.452 40.271 ;
    RECT 0.000 40.271 57.452 39.854 ;
    RECT 0.140 39.854 57.452 39.714 ;
    RECT 0.000 39.714 57.452 39.296 ;
    RECT 0.140 39.296 57.452 39.156 ;
    RECT 0.000 39.156 57.452 38.739 ;
    RECT 0.140 38.739 57.452 38.599 ;
    RECT 0.000 38.599 57.452 38.182 ;
    RECT 0.140 38.182 57.452 38.042 ;
    RECT 0.000 38.042 57.452 37.624 ;
    RECT 0.140 37.624 57.452 37.484 ;
    RECT 0.000 37.484 57.452 37.067 ;
    RECT 0.140 37.067 57.452 36.927 ;
    RECT 0.000 36.927 57.452 36.510 ;
    RECT 0.140 36.510 57.452 36.370 ;
    RECT 0.000 36.370 57.452 35.952 ;
    RECT 0.140 35.952 57.452 35.812 ;
    RECT 0.000 35.812 57.452 35.395 ;
    RECT 0.140 35.395 57.452 35.255 ;
    RECT 0.000 35.255 57.452 34.838 ;
    RECT 0.140 34.838 57.452 34.698 ;
    RECT 0.000 34.698 57.452 34.281 ;
    RECT 0.140 34.281 57.452 34.141 ;
    RECT 0.000 34.141 57.452 33.723 ;
    RECT 0.140 33.723 57.452 33.583 ;
    RECT 0.000 33.583 57.452 33.166 ;
    RECT 0.140 33.166 57.452 33.026 ;
    RECT 0.000 33.026 57.452 32.609 ;
    RECT 0.140 32.609 57.452 32.469 ;
    RECT 0.000 32.469 57.452 32.051 ;
    RECT 0.140 32.051 57.452 31.911 ;
    RECT 0.000 31.911 57.452 31.494 ;
    RECT 0.140 31.494 57.452 31.354 ;
    RECT 0.000 31.354 57.452 30.937 ;
    RECT 0.140 30.937 57.452 30.797 ;
    RECT 0.000 30.797 57.452 30.379 ;
    RECT 0.140 30.379 57.452 30.239 ;
    RECT 0.000 30.239 57.452 29.822 ;
    RECT 0.140 29.822 57.452 29.682 ;
    RECT 0.000 29.682 57.452 29.265 ;
    RECT 0.140 29.265 57.452 29.125 ;
    RECT 0.000 29.125 57.452 28.708 ;
    RECT 0.140 28.708 57.452 28.568 ;
    RECT 0.000 28.568 57.452 28.150 ;
    RECT 0.140 28.150 57.452 28.010 ;
    RECT 0.000 28.010 57.452 27.593 ;
    RECT 0.140 27.593 57.452 27.453 ;
    RECT 0.000 27.453 57.452 27.036 ;
    RECT 0.140 27.036 57.452 26.896 ;
    RECT 0.000 26.896 57.452 26.478 ;
    RECT 0.140 26.478 57.452 26.338 ;
    RECT 0.000 26.338 57.452 25.921 ;
    RECT 0.140 25.921 57.452 25.781 ;
    RECT 0.000 25.781 57.452 25.364 ;
    RECT 0.140 25.364 57.452 25.224 ;
    RECT 0.000 25.224 57.452 24.807 ;
    RECT 0.140 24.807 57.452 24.667 ;
    RECT 0.000 24.667 57.452 24.249 ;
    RECT 0.140 24.249 57.452 24.109 ;
    RECT 0.000 24.109 57.452 23.692 ;
    RECT 0.140 23.692 57.452 23.552 ;
    RECT 0.000 23.552 57.452 23.135 ;
    RECT 0.140 23.135 57.452 22.995 ;
    RECT 0.000 22.995 57.452 22.577 ;
    RECT 0.140 22.577 57.452 22.437 ;
    RECT 0.000 22.437 57.452 22.020 ;
    RECT 0.140 22.020 57.452 21.880 ;
    RECT 0.000 21.880 57.452 21.463 ;
    RECT 0.140 21.463 57.452 21.323 ;
    RECT 0.000 21.323 57.452 20.905 ;
    RECT 0.140 20.905 57.452 20.765 ;
    RECT 0.000 20.765 57.452 20.348 ;
    RECT 0.140 20.348 57.452 20.208 ;
    RECT 0.000 20.208 57.452 19.791 ;
    RECT 0.140 19.791 57.452 19.651 ;
    RECT 0.000 19.651 57.452 19.234 ;
    RECT 0.140 19.234 57.452 19.094 ;
    RECT 0.000 19.094 57.452 18.676 ;
    RECT 0.140 18.676 57.452 18.536 ;
    RECT 0.000 18.536 57.452 18.119 ;
    RECT 0.140 18.119 57.452 17.979 ;
    RECT 0.000 17.979 57.452 17.562 ;
    RECT 0.140 17.562 57.452 17.422 ;
    RECT 0.000 17.422 57.452 17.004 ;
    RECT 0.140 17.004 57.452 16.864 ;
    RECT 0.000 16.864 57.452 16.447 ;
    RECT 0.140 16.447 57.452 16.307 ;
    RECT 0.000 16.307 57.452 15.890 ;
    RECT 0.140 15.890 57.452 15.750 ;
    RECT 0.000 15.750 57.452 15.332 ;
    RECT 0.140 15.332 57.452 15.192 ;
    RECT 0.000 15.192 57.452 14.775 ;
    RECT 0.140 14.775 57.452 14.635 ;
    RECT 0.000 14.635 57.452 14.218 ;
    RECT 0.140 14.218 57.452 14.078 ;
    RECT 0.000 14.078 57.452 13.661 ;
    RECT 0.140 13.661 57.452 13.521 ;
    RECT 0.000 13.521 57.452 13.103 ;
    RECT 0.140 13.103 57.452 12.963 ;
    RECT 0.000 12.963 57.452 12.546 ;
    RECT 0.140 12.546 57.452 12.406 ;
    RECT 0.000 12.406 57.452 11.989 ;
    RECT 0.140 11.989 57.452 11.849 ;
    RECT 0.000 11.849 57.452 11.431 ;
    RECT 0.140 11.431 57.452 11.291 ;
    RECT 0.000 11.291 57.452 10.874 ;
    RECT 0.140 10.874 57.452 10.734 ;
    RECT 0.000 10.734 57.452 10.317 ;
    RECT 0.140 10.317 57.452 10.177 ;
    RECT 0.000 10.177 57.452 9.759 ;
    RECT 0.140 9.759 57.452 9.619 ;
    RECT 0.000 9.619 57.452 9.202 ;
    RECT 0.140 9.202 57.452 9.062 ;
    RECT 0.000 9.062 57.452 8.645 ;
    RECT 0.140 8.645 57.452 8.505 ;
    RECT 0.000 8.505 57.452 8.088 ;
    RECT 0.140 8.088 57.452 7.948 ;
    RECT 0.000 7.948 57.452 7.530 ;
    RECT 0.140 7.530 57.452 7.390 ;
    RECT 0.000 7.390 57.452 6.973 ;
    RECT 0.140 6.973 57.452 6.833 ;
    RECT 0.000 6.833 57.452 6.416 ;
    RECT 0.140 6.416 57.452 6.276 ;
    RECT 0.000 6.276 57.452 5.858 ;
    RECT 0.140 5.858 57.452 5.718 ;
    RECT 0.000 5.718 57.452 5.301 ;
    RECT 0.140 5.301 57.452 5.161 ;
    RECT 0.000 5.161 57.452 4.744 ;
    RECT 0.140 4.744 57.452 4.604 ;
    RECT 0.000 4.604 57.452 4.186 ;
    RECT 0.140 4.186 57.452 4.046 ;
    RECT 0.000 4.046 57.452 3.629 ;
    RECT 0.140 3.629 57.452 3.489 ;
    RECT 0.000 3.489 57.452 3.072 ;
    RECT 0.140 3.072 57.452 2.932 ;
    RECT 0.000 2.932 57.452 2.515 ;
    RECT 0.140 2.515 57.452 2.375 ;
    RECT 0.000 2.375 57.452 1.957 ;
    RECT 0.140 1.957 57.452 1.817 ;
    RECT 0.000 1.817 57.452 1.400 ;
    RECT 0.000 1.400 57.452 0.000 ;
    LAYER OVERLAP ;
    RECT 0 0 57.452 167.760 ;
    END
  END fakeram45_256x95

END LIBRARY
