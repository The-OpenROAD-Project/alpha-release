VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x15
  FOREIGN fakeram45_64x15 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 14.274 BY 41.681 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 40.141 0.140 40.281 ;
      LAYER metal2 ;
      RECT 0.000 40.141 0.140 40.281 ;
      LAYER metal3 ;
      RECT 0.000 40.141 0.140 40.281 ;
      LAYER metal4 ;
      RECT 0.000 40.141 0.140 40.281 ;
      END
    END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 39.421 0.140 39.561 ;
      LAYER metal2 ;
      RECT 0.000 39.421 0.140 39.561 ;
      LAYER metal3 ;
      RECT 0.000 39.421 0.140 39.561 ;
      LAYER metal4 ;
      RECT 0.000 39.421 0.140 39.561 ;
      END
    END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 38.701 0.140 38.841 ;
      LAYER metal2 ;
      RECT 0.000 38.701 0.140 38.841 ;
      LAYER metal3 ;
      RECT 0.000 38.701 0.140 38.841 ;
      LAYER metal4 ;
      RECT 0.000 38.701 0.140 38.841 ;
      END
    END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 37.981 0.140 38.121 ;
      LAYER metal2 ;
      RECT 0.000 37.981 0.140 38.121 ;
      LAYER metal3 ;
      RECT 0.000 37.981 0.140 38.121 ;
      LAYER metal4 ;
      RECT 0.000 37.981 0.140 38.121 ;
      END
    END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 37.261 0.140 37.401 ;
      LAYER metal2 ;
      RECT 0.000 37.261 0.140 37.401 ;
      LAYER metal3 ;
      RECT 0.000 37.261 0.140 37.401 ;
      LAYER metal4 ;
      RECT 0.000 37.261 0.140 37.401 ;
      END
    END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 36.541 0.140 36.681 ;
      LAYER metal2 ;
      RECT 0.000 36.541 0.140 36.681 ;
      LAYER metal3 ;
      RECT 0.000 36.541 0.140 36.681 ;
      LAYER metal4 ;
      RECT 0.000 36.541 0.140 36.681 ;
      END
    END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 35.821 0.140 35.961 ;
      LAYER metal2 ;
      RECT 0.000 35.821 0.140 35.961 ;
      LAYER metal3 ;
      RECT 0.000 35.821 0.140 35.961 ;
      LAYER metal4 ;
      RECT 0.000 35.821 0.140 35.961 ;
      END
    END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 35.101 0.140 35.241 ;
      LAYER metal2 ;
      RECT 0.000 35.101 0.140 35.241 ;
      LAYER metal3 ;
      RECT 0.000 35.101 0.140 35.241 ;
      LAYER metal4 ;
      RECT 0.000 35.101 0.140 35.241 ;
      END
    END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 34.381 0.140 34.521 ;
      LAYER metal2 ;
      RECT 0.000 34.381 0.140 34.521 ;
      LAYER metal3 ;
      RECT 0.000 34.381 0.140 34.521 ;
      LAYER metal4 ;
      RECT 0.000 34.381 0.140 34.521 ;
      END
    END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 33.661 0.140 33.801 ;
      LAYER metal2 ;
      RECT 0.000 33.661 0.140 33.801 ;
      LAYER metal3 ;
      RECT 0.000 33.661 0.140 33.801 ;
      LAYER metal4 ;
      RECT 0.000 33.661 0.140 33.801 ;
      END
    END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 32.941 0.140 33.081 ;
      LAYER metal2 ;
      RECT 0.000 32.941 0.140 33.081 ;
      LAYER metal3 ;
      RECT 0.000 32.941 0.140 33.081 ;
      LAYER metal4 ;
      RECT 0.000 32.941 0.140 33.081 ;
      END
    END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 32.221 0.140 32.361 ;
      LAYER metal2 ;
      RECT 0.000 32.221 0.140 32.361 ;
      LAYER metal3 ;
      RECT 0.000 32.221 0.140 32.361 ;
      LAYER metal4 ;
      RECT 0.000 32.221 0.140 32.361 ;
      END
    END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 31.501 0.140 31.641 ;
      LAYER metal2 ;
      RECT 0.000 31.501 0.140 31.641 ;
      LAYER metal3 ;
      RECT 0.000 31.501 0.140 31.641 ;
      LAYER metal4 ;
      RECT 0.000 31.501 0.140 31.641 ;
      END
    END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 30.781 0.140 30.921 ;
      LAYER metal2 ;
      RECT 0.000 30.781 0.140 30.921 ;
      LAYER metal3 ;
      RECT 0.000 30.781 0.140 30.921 ;
      LAYER metal4 ;
      RECT 0.000 30.781 0.140 30.921 ;
      END
    END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 30.061 0.140 30.201 ;
      LAYER metal2 ;
      RECT 0.000 30.061 0.140 30.201 ;
      LAYER metal3 ;
      RECT 0.000 30.061 0.140 30.201 ;
      LAYER metal4 ;
      RECT 0.000 30.061 0.140 30.201 ;
      END
    END w_mask_in[14]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 29.341 0.140 29.481 ;
      LAYER metal2 ;
      RECT 0.000 29.341 0.140 29.481 ;
      LAYER metal3 ;
      RECT 0.000 29.341 0.140 29.481 ;
      LAYER metal4 ;
      RECT 0.000 29.341 0.140 29.481 ;
      END
    END we_in
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 28.621 0.140 28.761 ;
      LAYER metal2 ;
      RECT 0.000 28.621 0.140 28.761 ;
      LAYER metal3 ;
      RECT 0.000 28.621 0.140 28.761 ;
      LAYER metal4 ;
      RECT 0.000 28.621 0.140 28.761 ;
      END
    END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 27.901 0.140 28.041 ;
      LAYER metal2 ;
      RECT 0.000 27.901 0.140 28.041 ;
      LAYER metal3 ;
      RECT 0.000 27.901 0.140 28.041 ;
      LAYER metal4 ;
      RECT 0.000 27.901 0.140 28.041 ;
      END
    END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 27.181 0.140 27.321 ;
      LAYER metal2 ;
      RECT 0.000 27.181 0.140 27.321 ;
      LAYER metal3 ;
      RECT 0.000 27.181 0.140 27.321 ;
      LAYER metal4 ;
      RECT 0.000 27.181 0.140 27.321 ;
      END
    END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 26.461 0.140 26.601 ;
      LAYER metal2 ;
      RECT 0.000 26.461 0.140 26.601 ;
      LAYER metal3 ;
      RECT 0.000 26.461 0.140 26.601 ;
      LAYER metal4 ;
      RECT 0.000 26.461 0.140 26.601 ;
      END
    END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 25.741 0.140 25.881 ;
      LAYER metal2 ;
      RECT 0.000 25.741 0.140 25.881 ;
      LAYER metal3 ;
      RECT 0.000 25.741 0.140 25.881 ;
      LAYER metal4 ;
      RECT 0.000 25.741 0.140 25.881 ;
      END
    END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 25.021 0.140 25.161 ;
      LAYER metal2 ;
      RECT 0.000 25.021 0.140 25.161 ;
      LAYER metal3 ;
      RECT 0.000 25.021 0.140 25.161 ;
      LAYER metal4 ;
      RECT 0.000 25.021 0.140 25.161 ;
      END
    END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 24.301 0.140 24.441 ;
      LAYER metal2 ;
      RECT 0.000 24.301 0.140 24.441 ;
      LAYER metal3 ;
      RECT 0.000 24.301 0.140 24.441 ;
      LAYER metal4 ;
      RECT 0.000 24.301 0.140 24.441 ;
      END
    END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 23.581 0.140 23.721 ;
      LAYER metal2 ;
      RECT 0.000 23.581 0.140 23.721 ;
      LAYER metal3 ;
      RECT 0.000 23.581 0.140 23.721 ;
      LAYER metal4 ;
      RECT 0.000 23.581 0.140 23.721 ;
      END
    END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 22.861 0.140 23.001 ;
      LAYER metal2 ;
      RECT 0.000 22.861 0.140 23.001 ;
      LAYER metal3 ;
      RECT 0.000 22.861 0.140 23.001 ;
      LAYER metal4 ;
      RECT 0.000 22.861 0.140 23.001 ;
      END
    END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 22.141 0.140 22.281 ;
      LAYER metal2 ;
      RECT 0.000 22.141 0.140 22.281 ;
      LAYER metal3 ;
      RECT 0.000 22.141 0.140 22.281 ;
      LAYER metal4 ;
      RECT 0.000 22.141 0.140 22.281 ;
      END
    END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 21.421 0.140 21.561 ;
      LAYER metal2 ;
      RECT 0.000 21.421 0.140 21.561 ;
      LAYER metal3 ;
      RECT 0.000 21.421 0.140 21.561 ;
      LAYER metal4 ;
      RECT 0.000 21.421 0.140 21.561 ;
      END
    END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 20.701 0.140 20.841 ;
      LAYER metal2 ;
      RECT 0.000 20.701 0.140 20.841 ;
      LAYER metal3 ;
      RECT 0.000 20.701 0.140 20.841 ;
      LAYER metal4 ;
      RECT 0.000 20.701 0.140 20.841 ;
      END
    END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 19.981 0.140 20.121 ;
      LAYER metal2 ;
      RECT 0.000 19.981 0.140 20.121 ;
      LAYER metal3 ;
      RECT 0.000 19.981 0.140 20.121 ;
      LAYER metal4 ;
      RECT 0.000 19.981 0.140 20.121 ;
      END
    END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 19.261 0.140 19.401 ;
      LAYER metal2 ;
      RECT 0.000 19.261 0.140 19.401 ;
      LAYER metal3 ;
      RECT 0.000 19.261 0.140 19.401 ;
      LAYER metal4 ;
      RECT 0.000 19.261 0.140 19.401 ;
      END
    END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 18.541 0.140 18.681 ;
      LAYER metal2 ;
      RECT 0.000 18.541 0.140 18.681 ;
      LAYER metal3 ;
      RECT 0.000 18.541 0.140 18.681 ;
      LAYER metal4 ;
      RECT 0.000 18.541 0.140 18.681 ;
      END
    END rd_out[14]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 17.820 0.140 17.960 ;
      LAYER metal2 ;
      RECT 0.000 17.820 0.140 17.960 ;
      LAYER metal3 ;
      RECT 0.000 17.820 0.140 17.960 ;
      LAYER metal4 ;
      RECT 0.000 17.820 0.140 17.960 ;
      END
    END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 17.100 0.140 17.240 ;
      LAYER metal2 ;
      RECT 0.000 17.100 0.140 17.240 ;
      LAYER metal3 ;
      RECT 0.000 17.100 0.140 17.240 ;
      LAYER metal4 ;
      RECT 0.000 17.100 0.140 17.240 ;
      END
    END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 16.380 0.140 16.520 ;
      LAYER metal2 ;
      RECT 0.000 16.380 0.140 16.520 ;
      LAYER metal3 ;
      RECT 0.000 16.380 0.140 16.520 ;
      LAYER metal4 ;
      RECT 0.000 16.380 0.140 16.520 ;
      END
    END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 15.660 0.140 15.800 ;
      LAYER metal2 ;
      RECT 0.000 15.660 0.140 15.800 ;
      LAYER metal3 ;
      RECT 0.000 15.660 0.140 15.800 ;
      LAYER metal4 ;
      RECT 0.000 15.660 0.140 15.800 ;
      END
    END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 14.940 0.140 15.080 ;
      LAYER metal2 ;
      RECT 0.000 14.940 0.140 15.080 ;
      LAYER metal3 ;
      RECT 0.000 14.940 0.140 15.080 ;
      LAYER metal4 ;
      RECT 0.000 14.940 0.140 15.080 ;
      END
    END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 14.220 0.140 14.360 ;
      LAYER metal2 ;
      RECT 0.000 14.220 0.140 14.360 ;
      LAYER metal3 ;
      RECT 0.000 14.220 0.140 14.360 ;
      LAYER metal4 ;
      RECT 0.000 14.220 0.140 14.360 ;
      END
    END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 13.500 0.140 13.640 ;
      LAYER metal2 ;
      RECT 0.000 13.500 0.140 13.640 ;
      LAYER metal3 ;
      RECT 0.000 13.500 0.140 13.640 ;
      LAYER metal4 ;
      RECT 0.000 13.500 0.140 13.640 ;
      END
    END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 12.780 0.140 12.920 ;
      LAYER metal2 ;
      RECT 0.000 12.780 0.140 12.920 ;
      LAYER metal3 ;
      RECT 0.000 12.780 0.140 12.920 ;
      LAYER metal4 ;
      RECT 0.000 12.780 0.140 12.920 ;
      END
    END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 12.060 0.140 12.200 ;
      LAYER metal2 ;
      RECT 0.000 12.060 0.140 12.200 ;
      LAYER metal3 ;
      RECT 0.000 12.060 0.140 12.200 ;
      LAYER metal4 ;
      RECT 0.000 12.060 0.140 12.200 ;
      END
    END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 11.340 0.140 11.480 ;
      LAYER metal2 ;
      RECT 0.000 11.340 0.140 11.480 ;
      LAYER metal3 ;
      RECT 0.000 11.340 0.140 11.480 ;
      LAYER metal4 ;
      RECT 0.000 11.340 0.140 11.480 ;
      END
    END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 10.620 0.140 10.760 ;
      LAYER metal2 ;
      RECT 0.000 10.620 0.140 10.760 ;
      LAYER metal3 ;
      RECT 0.000 10.620 0.140 10.760 ;
      LAYER metal4 ;
      RECT 0.000 10.620 0.140 10.760 ;
      END
    END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 9.900 0.140 10.040 ;
      LAYER metal2 ;
      RECT 0.000 9.900 0.140 10.040 ;
      LAYER metal3 ;
      RECT 0.000 9.900 0.140 10.040 ;
      LAYER metal4 ;
      RECT 0.000 9.900 0.140 10.040 ;
      END
    END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 9.180 0.140 9.320 ;
      LAYER metal2 ;
      RECT 0.000 9.180 0.140 9.320 ;
      LAYER metal3 ;
      RECT 0.000 9.180 0.140 9.320 ;
      LAYER metal4 ;
      RECT 0.000 9.180 0.140 9.320 ;
      END
    END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 8.460 0.140 8.600 ;
      LAYER metal2 ;
      RECT 0.000 8.460 0.140 8.600 ;
      LAYER metal3 ;
      RECT 0.000 8.460 0.140 8.600 ;
      LAYER metal4 ;
      RECT 0.000 8.460 0.140 8.600 ;
      END
    END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 7.740 0.140 7.880 ;
      LAYER metal2 ;
      RECT 0.000 7.740 0.140 7.880 ;
      LAYER metal3 ;
      RECT 0.000 7.740 0.140 7.880 ;
      LAYER metal4 ;
      RECT 0.000 7.740 0.140 7.880 ;
      END
    END wd_in[14]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 7.020 0.140 7.160 ;
      LAYER metal2 ;
      RECT 0.000 7.020 0.140 7.160 ;
      LAYER metal3 ;
      RECT 0.000 7.020 0.140 7.160 ;
      LAYER metal4 ;
      RECT 0.000 7.020 0.140 7.160 ;
      END
    END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 6.300 0.140 6.440 ;
      LAYER metal2 ;
      RECT 0.000 6.300 0.140 6.440 ;
      LAYER metal3 ;
      RECT 0.000 6.300 0.140 6.440 ;
      LAYER metal4 ;
      RECT 0.000 6.300 0.140 6.440 ;
      END
    END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 5.580 0.140 5.720 ;
      LAYER metal2 ;
      RECT 0.000 5.580 0.140 5.720 ;
      LAYER metal3 ;
      RECT 0.000 5.580 0.140 5.720 ;
      LAYER metal4 ;
      RECT 0.000 5.580 0.140 5.720 ;
      END
    END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 4.860 0.140 5.000 ;
      LAYER metal2 ;
      RECT 0.000 4.860 0.140 5.000 ;
      LAYER metal3 ;
      RECT 0.000 4.860 0.140 5.000 ;
      LAYER metal4 ;
      RECT 0.000 4.860 0.140 5.000 ;
      END
    END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 4.140 0.140 4.280 ;
      LAYER metal2 ;
      RECT 0.000 4.140 0.140 4.280 ;
      LAYER metal3 ;
      RECT 0.000 4.140 0.140 4.280 ;
      LAYER metal4 ;
      RECT 0.000 4.140 0.140 4.280 ;
      END
    END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 3.420 0.140 3.560 ;
      LAYER metal2 ;
      RECT 0.000 3.420 0.140 3.560 ;
      LAYER metal3 ;
      RECT 0.000 3.420 0.140 3.560 ;
      LAYER metal4 ;
      RECT 0.000 3.420 0.140 3.560 ;
      END
    END addr_in[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 2.700 0.140 2.840 ;
      LAYER metal2 ;
      RECT 0.000 2.700 0.140 2.840 ;
      LAYER metal3 ;
      RECT 0.000 2.700 0.140 2.840 ;
      LAYER metal4 ;
      RECT 0.000 2.700 0.140 2.840 ;
      END
    END clk
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
      RECT 0.000 1.980 0.140 2.120 ;
      LAYER metal2 ;
      RECT 0.000 1.980 0.140 2.120 ;
      LAYER metal3 ;
      RECT 0.000 1.980 0.140 2.120 ;
      LAYER metal4 ;
      RECT 0.000 1.980 0.140 2.120 ;
      END
    END ce_in
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.784 40.281 12.490 40.841 ;
      RECT 1.784 37.481 12.490 38.041 ;
      RECT 1.784 34.681 12.490 35.241 ;
      RECT 1.784 31.881 12.490 32.441 ;
      RECT 1.784 29.081 12.490 29.641 ;
      RECT 1.784 26.281 12.490 26.841 ;
      RECT 1.784 23.481 12.490 24.041 ;
      RECT 1.784 20.681 12.490 21.241 ;
      RECT 1.784 17.881 12.490 18.441 ;
      RECT 1.784 15.081 12.490 15.641 ;
      RECT 1.784 12.281 12.490 12.841 ;
      RECT 1.784 9.481 12.490 10.041 ;
      RECT 1.784 6.681 12.490 7.241 ;
      RECT 1.784 3.881 12.490 4.441 ;
      END
    END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 1.784 38.881 12.490 39.441 ;
      RECT 1.784 36.081 12.490 36.641 ;
      RECT 1.784 33.281 12.490 33.841 ;
      RECT 1.784 30.481 12.490 31.041 ;
      RECT 1.784 27.681 12.490 28.241 ;
      RECT 1.784 24.881 12.490 25.441 ;
      RECT 1.784 22.081 12.490 22.641 ;
      RECT 1.784 19.281 12.490 19.841 ;
      RECT 1.784 16.481 12.490 17.041 ;
      RECT 1.784 13.681 12.490 14.241 ;
      RECT 1.784 10.881 12.490 11.441 ;
      RECT 1.784 8.081 12.490 8.641 ;
      RECT 1.784 5.281 12.490 5.841 ;
      RECT 1.784 2.481 12.490 3.041 ;
      END
    END VDD
  OBS
    LAYER metal1 ;
    RECT 0.000 41.681 14.274 40.281 ;
    RECT 0.140 40.281 14.274 40.141 ;
    RECT 0.000 40.141 14.274 39.561 ;
    RECT 0.140 39.561 14.274 39.421 ;
    RECT 0.000 39.421 14.274 38.841 ;
    RECT 0.140 38.841 14.274 38.701 ;
    RECT 0.000 38.701 14.274 38.121 ;
    RECT 0.140 38.121 14.274 37.981 ;
    RECT 0.000 37.981 14.274 37.401 ;
    RECT 0.140 37.401 14.274 37.261 ;
    RECT 0.000 37.261 14.274 36.681 ;
    RECT 0.140 36.681 14.274 36.541 ;
    RECT 0.000 36.541 14.274 35.961 ;
    RECT 0.140 35.961 14.274 35.821 ;
    RECT 0.000 35.821 14.274 35.241 ;
    RECT 0.140 35.241 14.274 35.101 ;
    RECT 0.000 35.101 14.274 34.521 ;
    RECT 0.140 34.521 14.274 34.381 ;
    RECT 0.000 34.381 14.274 33.801 ;
    RECT 0.140 33.801 14.274 33.661 ;
    RECT 0.000 33.661 14.274 33.081 ;
    RECT 0.140 33.081 14.274 32.941 ;
    RECT 0.000 32.941 14.274 32.361 ;
    RECT 0.140 32.361 14.274 32.221 ;
    RECT 0.000 32.221 14.274 31.641 ;
    RECT 0.140 31.641 14.274 31.501 ;
    RECT 0.000 31.501 14.274 30.921 ;
    RECT 0.140 30.921 14.274 30.781 ;
    RECT 0.000 30.781 14.274 30.201 ;
    RECT 0.140 30.201 14.274 30.061 ;
    RECT 0.000 30.061 14.274 29.481 ;
    RECT 0.140 29.481 14.274 29.341 ;
    RECT 0.000 29.341 14.274 28.761 ;
    RECT 0.140 28.761 14.274 28.621 ;
    RECT 0.000 28.621 14.274 28.041 ;
    RECT 0.140 28.041 14.274 27.901 ;
    RECT 0.000 27.901 14.274 27.321 ;
    RECT 0.140 27.321 14.274 27.181 ;
    RECT 0.000 27.181 14.274 26.601 ;
    RECT 0.140 26.601 14.274 26.461 ;
    RECT 0.000 26.461 14.274 25.881 ;
    RECT 0.140 25.881 14.274 25.741 ;
    RECT 0.000 25.741 14.274 25.161 ;
    RECT 0.140 25.161 14.274 25.021 ;
    RECT 0.000 25.021 14.274 24.441 ;
    RECT 0.140 24.441 14.274 24.301 ;
    RECT 0.000 24.301 14.274 23.721 ;
    RECT 0.140 23.721 14.274 23.581 ;
    RECT 0.000 23.581 14.274 23.001 ;
    RECT 0.140 23.001 14.274 22.861 ;
    RECT 0.000 22.861 14.274 22.281 ;
    RECT 0.140 22.281 14.274 22.141 ;
    RECT 0.000 22.141 14.274 21.561 ;
    RECT 0.140 21.561 14.274 21.421 ;
    RECT 0.000 21.421 14.274 20.841 ;
    RECT 0.140 20.841 14.274 20.701 ;
    RECT 0.000 20.701 14.274 20.121 ;
    RECT 0.140 20.121 14.274 19.981 ;
    RECT 0.000 19.981 14.274 19.401 ;
    RECT 0.140 19.401 14.274 19.261 ;
    RECT 0.000 19.261 14.274 18.681 ;
    RECT 0.140 18.681 14.274 18.541 ;
    RECT 0.000 18.541 14.274 17.960 ;
    RECT 0.140 17.960 14.274 17.820 ;
    RECT 0.000 17.820 14.274 17.240 ;
    RECT 0.140 17.240 14.274 17.100 ;
    RECT 0.000 17.100 14.274 16.520 ;
    RECT 0.140 16.520 14.274 16.380 ;
    RECT 0.000 16.380 14.274 15.800 ;
    RECT 0.140 15.800 14.274 15.660 ;
    RECT 0.000 15.660 14.274 15.080 ;
    RECT 0.140 15.080 14.274 14.940 ;
    RECT 0.000 14.940 14.274 14.360 ;
    RECT 0.140 14.360 14.274 14.220 ;
    RECT 0.000 14.220 14.274 13.640 ;
    RECT 0.140 13.640 14.274 13.500 ;
    RECT 0.000 13.500 14.274 12.920 ;
    RECT 0.140 12.920 14.274 12.780 ;
    RECT 0.000 12.780 14.274 12.200 ;
    RECT 0.140 12.200 14.274 12.060 ;
    RECT 0.000 12.060 14.274 11.480 ;
    RECT 0.140 11.480 14.274 11.340 ;
    RECT 0.000 11.340 14.274 10.760 ;
    RECT 0.140 10.760 14.274 10.620 ;
    RECT 0.000 10.620 14.274 10.040 ;
    RECT 0.140 10.040 14.274 9.900 ;
    RECT 0.000 9.900 14.274 9.320 ;
    RECT 0.140 9.320 14.274 9.180 ;
    RECT 0.000 9.180 14.274 8.600 ;
    RECT 0.140 8.600 14.274 8.460 ;
    RECT 0.000 8.460 14.274 7.880 ;
    RECT 0.140 7.880 14.274 7.740 ;
    RECT 0.000 7.740 14.274 7.160 ;
    RECT 0.140 7.160 14.274 7.020 ;
    RECT 0.000 7.020 14.274 6.440 ;
    RECT 0.140 6.440 14.274 6.300 ;
    RECT 0.000 6.300 14.274 5.720 ;
    RECT 0.140 5.720 14.274 5.580 ;
    RECT 0.000 5.580 14.274 5.000 ;
    RECT 0.140 5.000 14.274 4.860 ;
    RECT 0.000 4.860 14.274 4.280 ;
    RECT 0.140 4.280 14.274 4.140 ;
    RECT 0.000 4.140 14.274 3.560 ;
    RECT 0.140 3.560 14.274 3.420 ;
    RECT 0.000 3.420 14.274 2.840 ;
    RECT 0.140 2.840 14.274 2.700 ;
    RECT 0.000 2.700 14.274 2.120 ;
    RECT 0.140 2.120 14.274 1.980 ;
    RECT 0.000 1.980 14.274 1.400 ;
    RECT 0.000 1.400 14.274 0.000 ;
    LAYER metal2 ;
    RECT 0.000 41.681 14.274 40.281 ;
    RECT 0.140 40.281 14.274 40.141 ;
    RECT 0.000 40.141 14.274 39.561 ;
    RECT 0.140 39.561 14.274 39.421 ;
    RECT 0.000 39.421 14.274 38.841 ;
    RECT 0.140 38.841 14.274 38.701 ;
    RECT 0.000 38.701 14.274 38.121 ;
    RECT 0.140 38.121 14.274 37.981 ;
    RECT 0.000 37.981 14.274 37.401 ;
    RECT 0.140 37.401 14.274 37.261 ;
    RECT 0.000 37.261 14.274 36.681 ;
    RECT 0.140 36.681 14.274 36.541 ;
    RECT 0.000 36.541 14.274 35.961 ;
    RECT 0.140 35.961 14.274 35.821 ;
    RECT 0.000 35.821 14.274 35.241 ;
    RECT 0.140 35.241 14.274 35.101 ;
    RECT 0.000 35.101 14.274 34.521 ;
    RECT 0.140 34.521 14.274 34.381 ;
    RECT 0.000 34.381 14.274 33.801 ;
    RECT 0.140 33.801 14.274 33.661 ;
    RECT 0.000 33.661 14.274 33.081 ;
    RECT 0.140 33.081 14.274 32.941 ;
    RECT 0.000 32.941 14.274 32.361 ;
    RECT 0.140 32.361 14.274 32.221 ;
    RECT 0.000 32.221 14.274 31.641 ;
    RECT 0.140 31.641 14.274 31.501 ;
    RECT 0.000 31.501 14.274 30.921 ;
    RECT 0.140 30.921 14.274 30.781 ;
    RECT 0.000 30.781 14.274 30.201 ;
    RECT 0.140 30.201 14.274 30.061 ;
    RECT 0.000 30.061 14.274 29.481 ;
    RECT 0.140 29.481 14.274 29.341 ;
    RECT 0.000 29.341 14.274 28.761 ;
    RECT 0.140 28.761 14.274 28.621 ;
    RECT 0.000 28.621 14.274 28.041 ;
    RECT 0.140 28.041 14.274 27.901 ;
    RECT 0.000 27.901 14.274 27.321 ;
    RECT 0.140 27.321 14.274 27.181 ;
    RECT 0.000 27.181 14.274 26.601 ;
    RECT 0.140 26.601 14.274 26.461 ;
    RECT 0.000 26.461 14.274 25.881 ;
    RECT 0.140 25.881 14.274 25.741 ;
    RECT 0.000 25.741 14.274 25.161 ;
    RECT 0.140 25.161 14.274 25.021 ;
    RECT 0.000 25.021 14.274 24.441 ;
    RECT 0.140 24.441 14.274 24.301 ;
    RECT 0.000 24.301 14.274 23.721 ;
    RECT 0.140 23.721 14.274 23.581 ;
    RECT 0.000 23.581 14.274 23.001 ;
    RECT 0.140 23.001 14.274 22.861 ;
    RECT 0.000 22.861 14.274 22.281 ;
    RECT 0.140 22.281 14.274 22.141 ;
    RECT 0.000 22.141 14.274 21.561 ;
    RECT 0.140 21.561 14.274 21.421 ;
    RECT 0.000 21.421 14.274 20.841 ;
    RECT 0.140 20.841 14.274 20.701 ;
    RECT 0.000 20.701 14.274 20.121 ;
    RECT 0.140 20.121 14.274 19.981 ;
    RECT 0.000 19.981 14.274 19.401 ;
    RECT 0.140 19.401 14.274 19.261 ;
    RECT 0.000 19.261 14.274 18.681 ;
    RECT 0.140 18.681 14.274 18.541 ;
    RECT 0.000 18.541 14.274 17.960 ;
    RECT 0.140 17.960 14.274 17.820 ;
    RECT 0.000 17.820 14.274 17.240 ;
    RECT 0.140 17.240 14.274 17.100 ;
    RECT 0.000 17.100 14.274 16.520 ;
    RECT 0.140 16.520 14.274 16.380 ;
    RECT 0.000 16.380 14.274 15.800 ;
    RECT 0.140 15.800 14.274 15.660 ;
    RECT 0.000 15.660 14.274 15.080 ;
    RECT 0.140 15.080 14.274 14.940 ;
    RECT 0.000 14.940 14.274 14.360 ;
    RECT 0.140 14.360 14.274 14.220 ;
    RECT 0.000 14.220 14.274 13.640 ;
    RECT 0.140 13.640 14.274 13.500 ;
    RECT 0.000 13.500 14.274 12.920 ;
    RECT 0.140 12.920 14.274 12.780 ;
    RECT 0.000 12.780 14.274 12.200 ;
    RECT 0.140 12.200 14.274 12.060 ;
    RECT 0.000 12.060 14.274 11.480 ;
    RECT 0.140 11.480 14.274 11.340 ;
    RECT 0.000 11.340 14.274 10.760 ;
    RECT 0.140 10.760 14.274 10.620 ;
    RECT 0.000 10.620 14.274 10.040 ;
    RECT 0.140 10.040 14.274 9.900 ;
    RECT 0.000 9.900 14.274 9.320 ;
    RECT 0.140 9.320 14.274 9.180 ;
    RECT 0.000 9.180 14.274 8.600 ;
    RECT 0.140 8.600 14.274 8.460 ;
    RECT 0.000 8.460 14.274 7.880 ;
    RECT 0.140 7.880 14.274 7.740 ;
    RECT 0.000 7.740 14.274 7.160 ;
    RECT 0.140 7.160 14.274 7.020 ;
    RECT 0.000 7.020 14.274 6.440 ;
    RECT 0.140 6.440 14.274 6.300 ;
    RECT 0.000 6.300 14.274 5.720 ;
    RECT 0.140 5.720 14.274 5.580 ;
    RECT 0.000 5.580 14.274 5.000 ;
    RECT 0.140 5.000 14.274 4.860 ;
    RECT 0.000 4.860 14.274 4.280 ;
    RECT 0.140 4.280 14.274 4.140 ;
    RECT 0.000 4.140 14.274 3.560 ;
    RECT 0.140 3.560 14.274 3.420 ;
    RECT 0.000 3.420 14.274 2.840 ;
    RECT 0.140 2.840 14.274 2.700 ;
    RECT 0.000 2.700 14.274 2.120 ;
    RECT 0.140 2.120 14.274 1.980 ;
    RECT 0.000 1.980 14.274 1.400 ;
    RECT 0.000 1.400 14.274 0.000 ;
    LAYER metal3 ;
    RECT 0.000 41.681 14.274 40.281 ;
    RECT 0.140 40.281 14.274 40.141 ;
    RECT 0.000 40.141 14.274 39.561 ;
    RECT 0.140 39.561 14.274 39.421 ;
    RECT 0.000 39.421 14.274 38.841 ;
    RECT 0.140 38.841 14.274 38.701 ;
    RECT 0.000 38.701 14.274 38.121 ;
    RECT 0.140 38.121 14.274 37.981 ;
    RECT 0.000 37.981 14.274 37.401 ;
    RECT 0.140 37.401 14.274 37.261 ;
    RECT 0.000 37.261 14.274 36.681 ;
    RECT 0.140 36.681 14.274 36.541 ;
    RECT 0.000 36.541 14.274 35.961 ;
    RECT 0.140 35.961 14.274 35.821 ;
    RECT 0.000 35.821 14.274 35.241 ;
    RECT 0.140 35.241 14.274 35.101 ;
    RECT 0.000 35.101 14.274 34.521 ;
    RECT 0.140 34.521 14.274 34.381 ;
    RECT 0.000 34.381 14.274 33.801 ;
    RECT 0.140 33.801 14.274 33.661 ;
    RECT 0.000 33.661 14.274 33.081 ;
    RECT 0.140 33.081 14.274 32.941 ;
    RECT 0.000 32.941 14.274 32.361 ;
    RECT 0.140 32.361 14.274 32.221 ;
    RECT 0.000 32.221 14.274 31.641 ;
    RECT 0.140 31.641 14.274 31.501 ;
    RECT 0.000 31.501 14.274 30.921 ;
    RECT 0.140 30.921 14.274 30.781 ;
    RECT 0.000 30.781 14.274 30.201 ;
    RECT 0.140 30.201 14.274 30.061 ;
    RECT 0.000 30.061 14.274 29.481 ;
    RECT 0.140 29.481 14.274 29.341 ;
    RECT 0.000 29.341 14.274 28.761 ;
    RECT 0.140 28.761 14.274 28.621 ;
    RECT 0.000 28.621 14.274 28.041 ;
    RECT 0.140 28.041 14.274 27.901 ;
    RECT 0.000 27.901 14.274 27.321 ;
    RECT 0.140 27.321 14.274 27.181 ;
    RECT 0.000 27.181 14.274 26.601 ;
    RECT 0.140 26.601 14.274 26.461 ;
    RECT 0.000 26.461 14.274 25.881 ;
    RECT 0.140 25.881 14.274 25.741 ;
    RECT 0.000 25.741 14.274 25.161 ;
    RECT 0.140 25.161 14.274 25.021 ;
    RECT 0.000 25.021 14.274 24.441 ;
    RECT 0.140 24.441 14.274 24.301 ;
    RECT 0.000 24.301 14.274 23.721 ;
    RECT 0.140 23.721 14.274 23.581 ;
    RECT 0.000 23.581 14.274 23.001 ;
    RECT 0.140 23.001 14.274 22.861 ;
    RECT 0.000 22.861 14.274 22.281 ;
    RECT 0.140 22.281 14.274 22.141 ;
    RECT 0.000 22.141 14.274 21.561 ;
    RECT 0.140 21.561 14.274 21.421 ;
    RECT 0.000 21.421 14.274 20.841 ;
    RECT 0.140 20.841 14.274 20.701 ;
    RECT 0.000 20.701 14.274 20.121 ;
    RECT 0.140 20.121 14.274 19.981 ;
    RECT 0.000 19.981 14.274 19.401 ;
    RECT 0.140 19.401 14.274 19.261 ;
    RECT 0.000 19.261 14.274 18.681 ;
    RECT 0.140 18.681 14.274 18.541 ;
    RECT 0.000 18.541 14.274 17.960 ;
    RECT 0.140 17.960 14.274 17.820 ;
    RECT 0.000 17.820 14.274 17.240 ;
    RECT 0.140 17.240 14.274 17.100 ;
    RECT 0.000 17.100 14.274 16.520 ;
    RECT 0.140 16.520 14.274 16.380 ;
    RECT 0.000 16.380 14.274 15.800 ;
    RECT 0.140 15.800 14.274 15.660 ;
    RECT 0.000 15.660 14.274 15.080 ;
    RECT 0.140 15.080 14.274 14.940 ;
    RECT 0.000 14.940 14.274 14.360 ;
    RECT 0.140 14.360 14.274 14.220 ;
    RECT 0.000 14.220 14.274 13.640 ;
    RECT 0.140 13.640 14.274 13.500 ;
    RECT 0.000 13.500 14.274 12.920 ;
    RECT 0.140 12.920 14.274 12.780 ;
    RECT 0.000 12.780 14.274 12.200 ;
    RECT 0.140 12.200 14.274 12.060 ;
    RECT 0.000 12.060 14.274 11.480 ;
    RECT 0.140 11.480 14.274 11.340 ;
    RECT 0.000 11.340 14.274 10.760 ;
    RECT 0.140 10.760 14.274 10.620 ;
    RECT 0.000 10.620 14.274 10.040 ;
    RECT 0.140 10.040 14.274 9.900 ;
    RECT 0.000 9.900 14.274 9.320 ;
    RECT 0.140 9.320 14.274 9.180 ;
    RECT 0.000 9.180 14.274 8.600 ;
    RECT 0.140 8.600 14.274 8.460 ;
    RECT 0.000 8.460 14.274 7.880 ;
    RECT 0.140 7.880 14.274 7.740 ;
    RECT 0.000 7.740 14.274 7.160 ;
    RECT 0.140 7.160 14.274 7.020 ;
    RECT 0.000 7.020 14.274 6.440 ;
    RECT 0.140 6.440 14.274 6.300 ;
    RECT 0.000 6.300 14.274 5.720 ;
    RECT 0.140 5.720 14.274 5.580 ;
    RECT 0.000 5.580 14.274 5.000 ;
    RECT 0.140 5.000 14.274 4.860 ;
    RECT 0.000 4.860 14.274 4.280 ;
    RECT 0.140 4.280 14.274 4.140 ;
    RECT 0.000 4.140 14.274 3.560 ;
    RECT 0.140 3.560 14.274 3.420 ;
    RECT 0.000 3.420 14.274 2.840 ;
    RECT 0.140 2.840 14.274 2.700 ;
    RECT 0.000 2.700 14.274 2.120 ;
    RECT 0.140 2.120 14.274 1.980 ;
    RECT 0.000 1.980 14.274 1.400 ;
    RECT 0.000 1.400 14.274 0.000 ;
    LAYER OVERLAP ;
    RECT 0 0 14.274 41.681 ;
    END
  END fakeram45_64x15

END LIBRARY
